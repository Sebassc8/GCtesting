
module aes_11cc ( clk, rst, g_init, e_init, o );
  input [127:0] g_init;
  input [127:0] e_init;
  output [127:0] o;
  input clk, rst;
  wire   N5, N6, N7, n7, \e/n291 , \e/n290 , \e/n289 , \e/n288 , \e/n287 ,
         \e/n286 , \e/n285 , \e/n284 , \e/n283 , \e/n282 , \e/n281 , \e/n280 ,
         \e/n279 , \e/n278 , \e/n277 , \e/n276 , \e/n275 , \e/n274 , \e/n273 ,
         \e/n272 , \e/n271 , \e/n270 , \e/n269 , \e/n268 , \e/n267 , \e/n266 ,
         \e/n265 , \e/n264 , \e/n263 , \e/n262 , \e/n261 , \e/n260 , \e/n259 ,
         \e/n258 , \e/n257 , \e/n256 , \e/n255 , \e/n254 , \e/n253 , \e/n252 ,
         \e/n251 , \e/n250 , \e/n249 , \e/n248 , \e/n247 , \e/n246 , \e/n245 ,
         \e/n244 , \e/n243 , \e/n242 , \e/n241 , \e/n240 , \e/n239 , \e/n238 ,
         \e/n237 , \e/n236 , \e/n235 , \e/n234 , \e/n233 , \e/n232 , \e/n231 ,
         \e/n230 , \e/n229 , \e/n228 , \e/n227 , \e/n226 , \e/n225 , \e/n224 ,
         \e/n223 , \e/n222 , \e/n221 , \e/n220 , \e/n219 , \e/n218 , \e/n217 ,
         \e/n216 , \e/n215 , \e/n214 , \e/n213 , \e/n212 , \e/n211 , \e/n210 ,
         \e/n209 , \e/n208 , \e/n207 , \e/n206 , \e/n205 , \e/n204 , \e/n203 ,
         \e/n202 , \e/n201 , \e/n200 , \e/n199 , \e/n198 , \e/n197 , \e/n196 ,
         \e/n195 , \e/n194 , \e/n193 , \e/n192 , \e/n191 , \e/n190 , \e/n189 ,
         \e/n188 , \e/n187 , \e/n186 , \e/n185 , \e/n184 , \e/n183 , \e/n182 ,
         \e/n181 , \e/n180 , \e/n178 , \e/n177 , \e/n176 , \e/n175 , \e/n174 ,
         \e/n173 , \e/n172 , \e/n171 , \e/n170 , \e/n169 , \e/n168 , \e/n167 ,
         \e/n166 , \e/n165 , \e/n164 , \e/n163 , \e/n162 , \e/n161 , \e/n160 ,
         \e/n159 , \e/n158 , \e/n157 , \e/n156 , \e/n155 , \e/n154 , \e/n153 ,
         \e/n152 , \e/n151 , \e/n150 , \e/n149 , \e/n148 , \e/n147 , \e/n98 ,
         \e/n97 , \e/n96 , \e/n95 , \e/n94 , \e/n93 , \e/n92 , \e/n91 ,
         \e/n90 , \e/n89 , \e/n88 , \e/n87 , \e/n86 , \e/n85 , \e/n84 ,
         \e/n83 , \e/n82 , \e/n81 , \e/n80 , \e/n79 , \e/n78 , \e/n77 ,
         \e/n76 , \e/n75 , \e/n74 , \e/n66 , \e/n58 , \e/n50 , \e/Q[7] ,
         \e/Q[4] , \e/Q[3] , \e/Q[2] , \e/t[10] , \e/t[11] , \e/t[12] ,
         \e/t[15] , \e/t[18] , \e/t[19] , \e/t[20] , \e/t[23] , \e/t[26] ,
         \e/t[27] , \e/t[28] , \e/t[31] , \e/w[3][0] , \e/w[3][1] ,
         \e/w[3][2] , \e/w[3][3] , \e/w[3][4] , \e/w[3][5] , \e/w[3][6] ,
         \e/w[3][7] , \e/w[3][8] , \e/w[3][9] , \e/w[3][10] , \e/w[3][11] ,
         \e/w[3][12] , \e/w[3][13] , \e/w[3][14] , \e/w[3][15] , \e/w[3][16] ,
         \e/w[3][17] , \e/w[3][18] , \e/w[3][19] , \e/w[3][20] , \e/w[3][21] ,
         \e/w[3][22] , \e/w[3][23] , \e/w[3][24] , \e/w[3][25] , \e/w[3][26] ,
         \e/w[3][27] , \e/w[3][28] , \e/w[3][29] , \e/w[3][30] , \e/w[3][31] ,
         \b/SBOX[0].sbox/n91 , \b/SBOX[0].sbox/n90 , \b/SBOX[0].sbox/n89 ,
         \b/SBOX[0].sbox/n88 , \b/SBOX[0].sbox/n87 , \b/SBOX[0].sbox/n86 ,
         \b/SBOX[0].sbox/n85 , \b/SBOX[0].sbox/n84 , \b/SBOX[0].sbox/n83 ,
         \b/SBOX[0].sbox/n82 , \b/SBOX[0].sbox/n81 , \b/SBOX[0].sbox/n80 ,
         \b/SBOX[0].sbox/n79 , \b/SBOX[0].sbox/n78 , \b/SBOX[0].sbox/n77 ,
         \b/SBOX[0].sbox/n76 , \b/SBOX[0].sbox/n75 , \b/SBOX[0].sbox/n74 ,
         \b/SBOX[0].sbox/n73 , \b/SBOX[0].sbox/n72 , \b/SBOX[0].sbox/n71 ,
         \b/SBOX[0].sbox/n70 , \b/SBOX[0].sbox/n69 , \b/SBOX[0].sbox/n68 ,
         \b/SBOX[0].sbox/n67 , \b/SBOX[0].sbox/n66 , \b/SBOX[0].sbox/n65 ,
         \b/SBOX[0].sbox/n64 , \b/SBOX[0].sbox/n63 , \b/SBOX[0].sbox/n62 ,
         \b/SBOX[0].sbox/n61 , \b/SBOX[0].sbox/n60 , \b/SBOX[0].sbox/n59 ,
         \b/SBOX[0].sbox/n58 , \b/SBOX[0].sbox/n57 , \b/SBOX[0].sbox/n56 ,
         \b/SBOX[0].sbox/n55 , \b/SBOX[0].sbox/n54 , \b/SBOX[0].sbox/n53 ,
         \b/SBOX[0].sbox/n52 , \b/SBOX[0].sbox/n51 , \b/SBOX[0].sbox/n50 ,
         \b/SBOX[0].sbox/n49 , \b/SBOX[0].sbox/n48 , \b/SBOX[0].sbox/n47 ,
         \b/SBOX[0].sbox/n46 , \b/SBOX[0].sbox/n45 , \b/SBOX[0].sbox/n44 ,
         \b/SBOX[0].sbox/n43 , \b/SBOX[0].sbox/n42 , \b/SBOX[0].sbox/n41 ,
         \b/SBOX[0].sbox/n40 , \b/SBOX[0].sbox/n39 , \b/SBOX[0].sbox/n38 ,
         \b/SBOX[0].sbox/n37 , \b/SBOX[0].sbox/n36 , \b/SBOX[0].sbox/n35 ,
         \b/SBOX[0].sbox/n34 , \b/SBOX[0].sbox/n33 , \b/SBOX[0].sbox/n32 ,
         \b/SBOX[0].sbox/n31 , \b/SBOX[0].sbox/n30 , \b/SBOX[0].sbox/n29 ,
         \b/SBOX[0].sbox/n28 , \b/SBOX[0].sbox/n27 , \b/SBOX[0].sbox/n26 ,
         \b/SBOX[0].sbox/n25 , \b/SBOX[0].sbox/n24 , \b/SBOX[0].sbox/n23 ,
         \b/SBOX[0].sbox/n22 , \b/SBOX[0].sbox/n21 , \b/SBOX[0].sbox/n20 ,
         \b/SBOX[0].sbox/n19 , \b/SBOX[0].sbox/n18 , \b/SBOX[0].sbox/n17 ,
         \b/SBOX[0].sbox/n16 , \b/SBOX[0].sbox/n15 , \b/SBOX[0].sbox/n14 ,
         \b/SBOX[0].sbox/n13 , \b/SBOX[0].sbox/n12 , \b/SBOX[0].sbox/n11 ,
         \b/SBOX[0].sbox/z[0] , \b/SBOX[0].sbox/z[1] , \b/SBOX[0].sbox/z[2] ,
         \b/SBOX[0].sbox/z[3] , \b/SBOX[0].sbox/z[4] , \b/SBOX[0].sbox/z[5] ,
         \b/SBOX[0].sbox/z[6] , \b/SBOX[0].sbox/z[7] , \b/SBOX[0].sbox/z[8] ,
         \b/SBOX[0].sbox/z[9] , \b/SBOX[0].sbox/z[10] , \b/SBOX[0].sbox/z[11] ,
         \b/SBOX[0].sbox/z[12] , \b/SBOX[0].sbox/z[13] ,
         \b/SBOX[0].sbox/z[14] , \b/SBOX[0].sbox/z[15] ,
         \b/SBOX[0].sbox/z[16] , \b/SBOX[0].sbox/z[17] , \b/SBOX[0].sbox/t[2] ,
         \b/SBOX[0].sbox/t[3] , \b/SBOX[0].sbox/t[5] , \b/SBOX[0].sbox/t[7] ,
         \b/SBOX[0].sbox/t[8] , \b/SBOX[0].sbox/t[10] , \b/SBOX[0].sbox/t[12] ,
         \b/SBOX[0].sbox/t[13] , \b/SBOX[0].sbox/t[15] ,
         \b/SBOX[0].sbox/t[21] , \b/SBOX[0].sbox/t[23] ,
         \b/SBOX[0].sbox/t[24] , \b/SBOX[0].sbox/t[25] ,
         \b/SBOX[0].sbox/t[26] , \b/SBOX[0].sbox/t[27] ,
         \b/SBOX[0].sbox/t[28] , \b/SBOX[0].sbox/t[29] ,
         \b/SBOX[0].sbox/t[30] , \b/SBOX[0].sbox/t[31] ,
         \b/SBOX[0].sbox/t[32] , \b/SBOX[0].sbox/t[33] ,
         \b/SBOX[0].sbox/t[36] , \b/SBOX[0].sbox/t[37] ,
         \b/SBOX[0].sbox/t[38] , \b/SBOX[0].sbox/t[39] ,
         \b/SBOX[0].sbox/t[40] , \b/SBOX[0].sbox/t[41] ,
         \b/SBOX[0].sbox/t[42] , \b/SBOX[0].sbox/t[43] ,
         \b/SBOX[0].sbox/t[44] , \b/SBOX[0].sbox/t[45] , \b/SBOX[0].sbox/y[1] ,
         \b/SBOX[0].sbox/y[2] , \b/SBOX[0].sbox/y[3] , \b/SBOX[0].sbox/y[4] ,
         \b/SBOX[0].sbox/y[5] , \b/SBOX[0].sbox/y[6] , \b/SBOX[0].sbox/y[7] ,
         \b/SBOX[0].sbox/y[10] , \b/SBOX[0].sbox/y[11] ,
         \b/SBOX[0].sbox/y[12] , \b/SBOX[0].sbox/y[15] ,
         \b/SBOX[0].sbox/y[16] , \b/SBOX[0].sbox/y[17] ,
         \e/a/SBOX[15].sbox/z[0] , \e/a/SBOX[15].sbox/z[1] ,
         \e/a/SBOX[15].sbox/z[2] , \e/a/SBOX[15].sbox/z[3] ,
         \e/a/SBOX[15].sbox/z[4] , \e/a/SBOX[15].sbox/z[5] ,
         \e/a/SBOX[15].sbox/z[6] , \e/a/SBOX[15].sbox/z[7] ,
         \e/a/SBOX[15].sbox/z[8] , \e/a/SBOX[15].sbox/z[9] ,
         \e/a/SBOX[15].sbox/z[10] , \e/a/SBOX[15].sbox/z[11] ,
         \e/a/SBOX[15].sbox/z[12] , \e/a/SBOX[15].sbox/z[13] ,
         \e/a/SBOX[15].sbox/z[14] , \e/a/SBOX[15].sbox/z[15] ,
         \e/a/SBOX[15].sbox/z[16] , \e/a/SBOX[15].sbox/z[17] ,
         \e/a/SBOX[15].sbox/t[2] , \e/a/SBOX[15].sbox/t[3] ,
         \e/a/SBOX[15].sbox/t[5] , \e/a/SBOX[15].sbox/t[7] ,
         \e/a/SBOX[15].sbox/t[8] , \e/a/SBOX[15].sbox/t[10] ,
         \e/a/SBOX[15].sbox/t[12] , \e/a/SBOX[15].sbox/t[13] ,
         \e/a/SBOX[15].sbox/t[15] , \e/a/SBOX[15].sbox/t[21] ,
         \e/a/SBOX[15].sbox/t[23] , \e/a/SBOX[15].sbox/t[24] ,
         \e/a/SBOX[15].sbox/t[25] , \e/a/SBOX[15].sbox/t[26] ,
         \e/a/SBOX[15].sbox/t[27] , \e/a/SBOX[15].sbox/t[28] ,
         \e/a/SBOX[15].sbox/t[29] , \e/a/SBOX[15].sbox/t[30] ,
         \e/a/SBOX[15].sbox/t[31] , \e/a/SBOX[15].sbox/t[32] ,
         \e/a/SBOX[15].sbox/t[33] , \e/a/SBOX[15].sbox/t[36] ,
         \e/a/SBOX[15].sbox/t[37] , \e/a/SBOX[15].sbox/t[38] ,
         \e/a/SBOX[15].sbox/t[39] , \e/a/SBOX[15].sbox/t[40] ,
         \e/a/SBOX[15].sbox/t[41] , \e/a/SBOX[15].sbox/t[42] ,
         \e/a/SBOX[15].sbox/t[43] , \e/a/SBOX[15].sbox/t[44] ,
         \e/a/SBOX[15].sbox/t[45] , \e/a/SBOX[15].sbox/y[1] ,
         \e/a/SBOX[15].sbox/y[2] , \e/a/SBOX[15].sbox/y[3] ,
         \e/a/SBOX[15].sbox/y[4] , \e/a/SBOX[15].sbox/y[5] ,
         \e/a/SBOX[15].sbox/y[6] , \e/a/SBOX[15].sbox/y[7] ,
         \e/a/SBOX[15].sbox/y[10] , \e/a/SBOX[15].sbox/y[11] ,
         \e/a/SBOX[15].sbox/y[12] , \e/a/SBOX[15].sbox/y[15] ,
         \e/a/SBOX[15].sbox/y[16] , \e/a/SBOX[15].sbox/y[17] ,
         \e/a/SBOX[14].sbox/z[0] , \e/a/SBOX[14].sbox/z[1] ,
         \e/a/SBOX[14].sbox/z[2] , \e/a/SBOX[14].sbox/z[3] ,
         \e/a/SBOX[14].sbox/z[4] , \e/a/SBOX[14].sbox/z[5] ,
         \e/a/SBOX[14].sbox/z[6] , \e/a/SBOX[14].sbox/z[7] ,
         \e/a/SBOX[14].sbox/z[8] , \e/a/SBOX[14].sbox/z[9] ,
         \e/a/SBOX[14].sbox/z[10] , \e/a/SBOX[14].sbox/z[11] ,
         \e/a/SBOX[14].sbox/z[12] , \e/a/SBOX[14].sbox/z[13] ,
         \e/a/SBOX[14].sbox/z[14] , \e/a/SBOX[14].sbox/z[15] ,
         \e/a/SBOX[14].sbox/z[16] , \e/a/SBOX[14].sbox/z[17] ,
         \e/a/SBOX[14].sbox/t[2] , \e/a/SBOX[14].sbox/t[3] ,
         \e/a/SBOX[14].sbox/t[5] , \e/a/SBOX[14].sbox/t[7] ,
         \e/a/SBOX[14].sbox/t[8] , \e/a/SBOX[14].sbox/t[10] ,
         \e/a/SBOX[14].sbox/t[12] , \e/a/SBOX[14].sbox/t[13] ,
         \e/a/SBOX[14].sbox/t[15] , \e/a/SBOX[14].sbox/t[21] ,
         \e/a/SBOX[14].sbox/t[23] , \e/a/SBOX[14].sbox/t[24] ,
         \e/a/SBOX[14].sbox/t[25] , \e/a/SBOX[14].sbox/t[26] ,
         \e/a/SBOX[14].sbox/t[27] , \e/a/SBOX[14].sbox/t[28] ,
         \e/a/SBOX[14].sbox/t[29] , \e/a/SBOX[14].sbox/t[30] ,
         \e/a/SBOX[14].sbox/t[31] , \e/a/SBOX[14].sbox/t[32] ,
         \e/a/SBOX[14].sbox/t[33] , \e/a/SBOX[14].sbox/t[36] ,
         \e/a/SBOX[14].sbox/t[37] , \e/a/SBOX[14].sbox/t[38] ,
         \e/a/SBOX[14].sbox/t[39] , \e/a/SBOX[14].sbox/t[40] ,
         \e/a/SBOX[14].sbox/t[41] , \e/a/SBOX[14].sbox/t[42] ,
         \e/a/SBOX[14].sbox/t[43] , \e/a/SBOX[14].sbox/t[44] ,
         \e/a/SBOX[14].sbox/t[45] , \e/a/SBOX[14].sbox/y[1] ,
         \e/a/SBOX[14].sbox/y[2] , \e/a/SBOX[14].sbox/y[3] ,
         \e/a/SBOX[14].sbox/y[4] , \e/a/SBOX[14].sbox/y[5] ,
         \e/a/SBOX[14].sbox/y[6] , \e/a/SBOX[14].sbox/y[7] ,
         \e/a/SBOX[14].sbox/y[10] , \e/a/SBOX[14].sbox/y[11] ,
         \e/a/SBOX[14].sbox/y[12] , \e/a/SBOX[14].sbox/y[15] ,
         \e/a/SBOX[14].sbox/y[16] , \e/a/SBOX[14].sbox/y[17] ,
         \e/a/SBOX[13].sbox/z[0] , \e/a/SBOX[13].sbox/z[1] ,
         \e/a/SBOX[13].sbox/z[2] , \e/a/SBOX[13].sbox/z[3] ,
         \e/a/SBOX[13].sbox/z[4] , \e/a/SBOX[13].sbox/z[5] ,
         \e/a/SBOX[13].sbox/z[6] , \e/a/SBOX[13].sbox/z[7] ,
         \e/a/SBOX[13].sbox/z[8] , \e/a/SBOX[13].sbox/z[9] ,
         \e/a/SBOX[13].sbox/z[10] , \e/a/SBOX[13].sbox/z[11] ,
         \e/a/SBOX[13].sbox/z[12] , \e/a/SBOX[13].sbox/z[13] ,
         \e/a/SBOX[13].sbox/z[14] , \e/a/SBOX[13].sbox/z[15] ,
         \e/a/SBOX[13].sbox/z[16] , \e/a/SBOX[13].sbox/z[17] ,
         \e/a/SBOX[13].sbox/t[2] , \e/a/SBOX[13].sbox/t[3] ,
         \e/a/SBOX[13].sbox/t[5] , \e/a/SBOX[13].sbox/t[7] ,
         \e/a/SBOX[13].sbox/t[8] , \e/a/SBOX[13].sbox/t[10] ,
         \e/a/SBOX[13].sbox/t[12] , \e/a/SBOX[13].sbox/t[13] ,
         \e/a/SBOX[13].sbox/t[15] , \e/a/SBOX[13].sbox/t[21] ,
         \e/a/SBOX[13].sbox/t[23] , \e/a/SBOX[13].sbox/t[24] ,
         \e/a/SBOX[13].sbox/t[25] , \e/a/SBOX[13].sbox/t[26] ,
         \e/a/SBOX[13].sbox/t[27] , \e/a/SBOX[13].sbox/t[28] ,
         \e/a/SBOX[13].sbox/t[29] , \e/a/SBOX[13].sbox/t[30] ,
         \e/a/SBOX[13].sbox/t[31] , \e/a/SBOX[13].sbox/t[32] ,
         \e/a/SBOX[13].sbox/t[33] , \e/a/SBOX[13].sbox/t[36] ,
         \e/a/SBOX[13].sbox/t[37] , \e/a/SBOX[13].sbox/t[38] ,
         \e/a/SBOX[13].sbox/t[39] , \e/a/SBOX[13].sbox/t[40] ,
         \e/a/SBOX[13].sbox/t[41] , \e/a/SBOX[13].sbox/t[42] ,
         \e/a/SBOX[13].sbox/t[43] , \e/a/SBOX[13].sbox/t[44] ,
         \e/a/SBOX[13].sbox/t[45] , \e/a/SBOX[13].sbox/y[1] ,
         \e/a/SBOX[13].sbox/y[2] , \e/a/SBOX[13].sbox/y[3] ,
         \e/a/SBOX[13].sbox/y[4] , \e/a/SBOX[13].sbox/y[5] ,
         \e/a/SBOX[13].sbox/y[6] , \e/a/SBOX[13].sbox/y[7] ,
         \e/a/SBOX[13].sbox/y[10] , \e/a/SBOX[13].sbox/y[11] ,
         \e/a/SBOX[13].sbox/y[12] , \e/a/SBOX[13].sbox/y[15] ,
         \e/a/SBOX[13].sbox/y[16] , \e/a/SBOX[13].sbox/y[17] ,
         \e/a/SBOX[12].sbox/z[0] , \e/a/SBOX[12].sbox/z[1] ,
         \e/a/SBOX[12].sbox/z[2] , \e/a/SBOX[12].sbox/z[3] ,
         \e/a/SBOX[12].sbox/z[4] , \e/a/SBOX[12].sbox/z[5] ,
         \e/a/SBOX[12].sbox/z[6] , \e/a/SBOX[12].sbox/z[7] ,
         \e/a/SBOX[12].sbox/z[8] , \e/a/SBOX[12].sbox/z[9] ,
         \e/a/SBOX[12].sbox/z[10] , \e/a/SBOX[12].sbox/z[11] ,
         \e/a/SBOX[12].sbox/z[12] , \e/a/SBOX[12].sbox/z[13] ,
         \e/a/SBOX[12].sbox/z[14] , \e/a/SBOX[12].sbox/z[15] ,
         \e/a/SBOX[12].sbox/z[16] , \e/a/SBOX[12].sbox/z[17] ,
         \e/a/SBOX[12].sbox/t[2] , \e/a/SBOX[12].sbox/t[3] ,
         \e/a/SBOX[12].sbox/t[5] , \e/a/SBOX[12].sbox/t[7] ,
         \e/a/SBOX[12].sbox/t[8] , \e/a/SBOX[12].sbox/t[10] ,
         \e/a/SBOX[12].sbox/t[12] , \e/a/SBOX[12].sbox/t[13] ,
         \e/a/SBOX[12].sbox/t[15] , \e/a/SBOX[12].sbox/t[21] ,
         \e/a/SBOX[12].sbox/t[23] , \e/a/SBOX[12].sbox/t[24] ,
         \e/a/SBOX[12].sbox/t[25] , \e/a/SBOX[12].sbox/t[26] ,
         \e/a/SBOX[12].sbox/t[27] , \e/a/SBOX[12].sbox/t[28] ,
         \e/a/SBOX[12].sbox/t[29] , \e/a/SBOX[12].sbox/t[30] ,
         \e/a/SBOX[12].sbox/t[31] , \e/a/SBOX[12].sbox/t[32] ,
         \e/a/SBOX[12].sbox/t[33] , \e/a/SBOX[12].sbox/t[36] ,
         \e/a/SBOX[12].sbox/t[37] , \e/a/SBOX[12].sbox/t[38] ,
         \e/a/SBOX[12].sbox/t[39] , \e/a/SBOX[12].sbox/t[40] ,
         \e/a/SBOX[12].sbox/t[41] , \e/a/SBOX[12].sbox/t[42] ,
         \e/a/SBOX[12].sbox/t[43] , \e/a/SBOX[12].sbox/t[44] ,
         \e/a/SBOX[12].sbox/t[45] , \e/a/SBOX[12].sbox/y[1] ,
         \e/a/SBOX[12].sbox/y[2] , \e/a/SBOX[12].sbox/y[3] ,
         \e/a/SBOX[12].sbox/y[4] , \e/a/SBOX[12].sbox/y[5] ,
         \e/a/SBOX[12].sbox/y[6] , \e/a/SBOX[12].sbox/y[7] ,
         \e/a/SBOX[12].sbox/y[10] , \e/a/SBOX[12].sbox/y[11] ,
         \e/a/SBOX[12].sbox/y[12] , \e/a/SBOX[12].sbox/y[15] ,
         \e/a/SBOX[12].sbox/y[16] , \e/a/SBOX[12].sbox/y[17] ,
         \b/SBOX[15].sbox/z[0] , \b/SBOX[15].sbox/z[1] ,
         \b/SBOX[15].sbox/z[2] , \b/SBOX[15].sbox/z[3] ,
         \b/SBOX[15].sbox/z[4] , \b/SBOX[15].sbox/z[5] ,
         \b/SBOX[15].sbox/z[6] , \b/SBOX[15].sbox/z[7] ,
         \b/SBOX[15].sbox/z[8] , \b/SBOX[15].sbox/z[9] ,
         \b/SBOX[15].sbox/z[10] , \b/SBOX[15].sbox/z[11] ,
         \b/SBOX[15].sbox/z[12] , \b/SBOX[15].sbox/z[13] ,
         \b/SBOX[15].sbox/z[14] , \b/SBOX[15].sbox/z[15] ,
         \b/SBOX[15].sbox/z[16] , \b/SBOX[15].sbox/z[17] ,
         \b/SBOX[15].sbox/t[2] , \b/SBOX[15].sbox/t[3] ,
         \b/SBOX[15].sbox/t[5] , \b/SBOX[15].sbox/t[7] ,
         \b/SBOX[15].sbox/t[8] , \b/SBOX[15].sbox/t[10] ,
         \b/SBOX[15].sbox/t[12] , \b/SBOX[15].sbox/t[13] ,
         \b/SBOX[15].sbox/t[15] , \b/SBOX[15].sbox/t[21] ,
         \b/SBOX[15].sbox/t[23] , \b/SBOX[15].sbox/t[24] ,
         \b/SBOX[15].sbox/t[25] , \b/SBOX[15].sbox/t[26] ,
         \b/SBOX[15].sbox/t[27] , \b/SBOX[15].sbox/t[28] ,
         \b/SBOX[15].sbox/t[29] , \b/SBOX[15].sbox/t[30] ,
         \b/SBOX[15].sbox/t[31] , \b/SBOX[15].sbox/t[32] ,
         \b/SBOX[15].sbox/t[33] , \b/SBOX[15].sbox/t[36] ,
         \b/SBOX[15].sbox/t[37] , \b/SBOX[15].sbox/t[38] ,
         \b/SBOX[15].sbox/t[39] , \b/SBOX[15].sbox/t[40] ,
         \b/SBOX[15].sbox/t[41] , \b/SBOX[15].sbox/t[42] ,
         \b/SBOX[15].sbox/t[43] , \b/SBOX[15].sbox/t[44] ,
         \b/SBOX[15].sbox/t[45] , \b/SBOX[15].sbox/y[1] ,
         \b/SBOX[15].sbox/y[2] , \b/SBOX[15].sbox/y[3] ,
         \b/SBOX[15].sbox/y[4] , \b/SBOX[15].sbox/y[5] ,
         \b/SBOX[15].sbox/y[6] , \b/SBOX[15].sbox/y[7] ,
         \b/SBOX[15].sbox/y[10] , \b/SBOX[15].sbox/y[11] ,
         \b/SBOX[15].sbox/y[12] , \b/SBOX[15].sbox/y[15] ,
         \b/SBOX[15].sbox/y[16] , \b/SBOX[15].sbox/y[17] ,
         \b/SBOX[14].sbox/z[0] , \b/SBOX[14].sbox/z[1] ,
         \b/SBOX[14].sbox/z[2] , \b/SBOX[14].sbox/z[3] ,
         \b/SBOX[14].sbox/z[4] , \b/SBOX[14].sbox/z[5] ,
         \b/SBOX[14].sbox/z[6] , \b/SBOX[14].sbox/z[7] ,
         \b/SBOX[14].sbox/z[8] , \b/SBOX[14].sbox/z[9] ,
         \b/SBOX[14].sbox/z[10] , \b/SBOX[14].sbox/z[11] ,
         \b/SBOX[14].sbox/z[12] , \b/SBOX[14].sbox/z[13] ,
         \b/SBOX[14].sbox/z[14] , \b/SBOX[14].sbox/z[15] ,
         \b/SBOX[14].sbox/z[16] , \b/SBOX[14].sbox/z[17] ,
         \b/SBOX[14].sbox/t[2] , \b/SBOX[14].sbox/t[3] ,
         \b/SBOX[14].sbox/t[5] , \b/SBOX[14].sbox/t[7] ,
         \b/SBOX[14].sbox/t[8] , \b/SBOX[14].sbox/t[10] ,
         \b/SBOX[14].sbox/t[12] , \b/SBOX[14].sbox/t[13] ,
         \b/SBOX[14].sbox/t[15] , \b/SBOX[14].sbox/t[21] ,
         \b/SBOX[14].sbox/t[23] , \b/SBOX[14].sbox/t[24] ,
         \b/SBOX[14].sbox/t[25] , \b/SBOX[14].sbox/t[26] ,
         \b/SBOX[14].sbox/t[27] , \b/SBOX[14].sbox/t[28] ,
         \b/SBOX[14].sbox/t[29] , \b/SBOX[14].sbox/t[30] ,
         \b/SBOX[14].sbox/t[31] , \b/SBOX[14].sbox/t[32] ,
         \b/SBOX[14].sbox/t[33] , \b/SBOX[14].sbox/t[36] ,
         \b/SBOX[14].sbox/t[37] , \b/SBOX[14].sbox/t[38] ,
         \b/SBOX[14].sbox/t[39] , \b/SBOX[14].sbox/t[40] ,
         \b/SBOX[14].sbox/t[41] , \b/SBOX[14].sbox/t[42] ,
         \b/SBOX[14].sbox/t[43] , \b/SBOX[14].sbox/t[44] ,
         \b/SBOX[14].sbox/t[45] , \b/SBOX[14].sbox/y[1] ,
         \b/SBOX[14].sbox/y[2] , \b/SBOX[14].sbox/y[3] ,
         \b/SBOX[14].sbox/y[4] , \b/SBOX[14].sbox/y[5] ,
         \b/SBOX[14].sbox/y[6] , \b/SBOX[14].sbox/y[7] ,
         \b/SBOX[14].sbox/y[10] , \b/SBOX[14].sbox/y[11] ,
         \b/SBOX[14].sbox/y[12] , \b/SBOX[14].sbox/y[15] ,
         \b/SBOX[14].sbox/y[16] , \b/SBOX[14].sbox/y[17] ,
         \b/SBOX[13].sbox/z[0] , \b/SBOX[13].sbox/z[1] ,
         \b/SBOX[13].sbox/z[2] , \b/SBOX[13].sbox/z[3] ,
         \b/SBOX[13].sbox/z[4] , \b/SBOX[13].sbox/z[5] ,
         \b/SBOX[13].sbox/z[6] , \b/SBOX[13].sbox/z[7] ,
         \b/SBOX[13].sbox/z[8] , \b/SBOX[13].sbox/z[9] ,
         \b/SBOX[13].sbox/z[10] , \b/SBOX[13].sbox/z[11] ,
         \b/SBOX[13].sbox/z[12] , \b/SBOX[13].sbox/z[13] ,
         \b/SBOX[13].sbox/z[14] , \b/SBOX[13].sbox/z[15] ,
         \b/SBOX[13].sbox/z[16] , \b/SBOX[13].sbox/z[17] ,
         \b/SBOX[13].sbox/t[2] , \b/SBOX[13].sbox/t[3] ,
         \b/SBOX[13].sbox/t[5] , \b/SBOX[13].sbox/t[7] ,
         \b/SBOX[13].sbox/t[8] , \b/SBOX[13].sbox/t[10] ,
         \b/SBOX[13].sbox/t[12] , \b/SBOX[13].sbox/t[13] ,
         \b/SBOX[13].sbox/t[15] , \b/SBOX[13].sbox/t[21] ,
         \b/SBOX[13].sbox/t[23] , \b/SBOX[13].sbox/t[24] ,
         \b/SBOX[13].sbox/t[25] , \b/SBOX[13].sbox/t[26] ,
         \b/SBOX[13].sbox/t[27] , \b/SBOX[13].sbox/t[28] ,
         \b/SBOX[13].sbox/t[29] , \b/SBOX[13].sbox/t[30] ,
         \b/SBOX[13].sbox/t[31] , \b/SBOX[13].sbox/t[32] ,
         \b/SBOX[13].sbox/t[33] , \b/SBOX[13].sbox/t[36] ,
         \b/SBOX[13].sbox/t[37] , \b/SBOX[13].sbox/t[38] ,
         \b/SBOX[13].sbox/t[39] , \b/SBOX[13].sbox/t[40] ,
         \b/SBOX[13].sbox/t[41] , \b/SBOX[13].sbox/t[42] ,
         \b/SBOX[13].sbox/t[43] , \b/SBOX[13].sbox/t[44] ,
         \b/SBOX[13].sbox/t[45] , \b/SBOX[13].sbox/y[1] ,
         \b/SBOX[13].sbox/y[2] , \b/SBOX[13].sbox/y[3] ,
         \b/SBOX[13].sbox/y[4] , \b/SBOX[13].sbox/y[5] ,
         \b/SBOX[13].sbox/y[6] , \b/SBOX[13].sbox/y[7] ,
         \b/SBOX[13].sbox/y[10] , \b/SBOX[13].sbox/y[11] ,
         \b/SBOX[13].sbox/y[12] , \b/SBOX[13].sbox/y[15] ,
         \b/SBOX[13].sbox/y[16] , \b/SBOX[13].sbox/y[17] ,
         \b/SBOX[12].sbox/z[0] , \b/SBOX[12].sbox/z[1] ,
         \b/SBOX[12].sbox/z[2] , \b/SBOX[12].sbox/z[3] ,
         \b/SBOX[12].sbox/z[4] , \b/SBOX[12].sbox/z[5] ,
         \b/SBOX[12].sbox/z[6] , \b/SBOX[12].sbox/z[7] ,
         \b/SBOX[12].sbox/z[8] , \b/SBOX[12].sbox/z[9] ,
         \b/SBOX[12].sbox/z[10] , \b/SBOX[12].sbox/z[11] ,
         \b/SBOX[12].sbox/z[12] , \b/SBOX[12].sbox/z[13] ,
         \b/SBOX[12].sbox/z[14] , \b/SBOX[12].sbox/z[15] ,
         \b/SBOX[12].sbox/z[16] , \b/SBOX[12].sbox/z[17] ,
         \b/SBOX[12].sbox/t[2] , \b/SBOX[12].sbox/t[3] ,
         \b/SBOX[12].sbox/t[5] , \b/SBOX[12].sbox/t[7] ,
         \b/SBOX[12].sbox/t[8] , \b/SBOX[12].sbox/t[10] ,
         \b/SBOX[12].sbox/t[12] , \b/SBOX[12].sbox/t[13] ,
         \b/SBOX[12].sbox/t[15] , \b/SBOX[12].sbox/t[21] ,
         \b/SBOX[12].sbox/t[23] , \b/SBOX[12].sbox/t[24] ,
         \b/SBOX[12].sbox/t[25] , \b/SBOX[12].sbox/t[26] ,
         \b/SBOX[12].sbox/t[27] , \b/SBOX[12].sbox/t[28] ,
         \b/SBOX[12].sbox/t[29] , \b/SBOX[12].sbox/t[30] ,
         \b/SBOX[12].sbox/t[31] , \b/SBOX[12].sbox/t[32] ,
         \b/SBOX[12].sbox/t[33] , \b/SBOX[12].sbox/t[36] ,
         \b/SBOX[12].sbox/t[37] , \b/SBOX[12].sbox/t[38] ,
         \b/SBOX[12].sbox/t[39] , \b/SBOX[12].sbox/t[40] ,
         \b/SBOX[12].sbox/t[41] , \b/SBOX[12].sbox/t[42] ,
         \b/SBOX[12].sbox/t[43] , \b/SBOX[12].sbox/t[44] ,
         \b/SBOX[12].sbox/t[45] , \b/SBOX[12].sbox/y[1] ,
         \b/SBOX[12].sbox/y[2] , \b/SBOX[12].sbox/y[3] ,
         \b/SBOX[12].sbox/y[4] , \b/SBOX[12].sbox/y[5] ,
         \b/SBOX[12].sbox/y[6] , \b/SBOX[12].sbox/y[7] ,
         \b/SBOX[12].sbox/y[10] , \b/SBOX[12].sbox/y[11] ,
         \b/SBOX[12].sbox/y[12] , \b/SBOX[12].sbox/y[15] ,
         \b/SBOX[12].sbox/y[16] , \b/SBOX[12].sbox/y[17] ,
         \b/SBOX[11].sbox/z[0] , \b/SBOX[11].sbox/z[1] ,
         \b/SBOX[11].sbox/z[2] , \b/SBOX[11].sbox/z[3] ,
         \b/SBOX[11].sbox/z[4] , \b/SBOX[11].sbox/z[5] ,
         \b/SBOX[11].sbox/z[6] , \b/SBOX[11].sbox/z[7] ,
         \b/SBOX[11].sbox/z[8] , \b/SBOX[11].sbox/z[9] ,
         \b/SBOX[11].sbox/z[10] , \b/SBOX[11].sbox/z[11] ,
         \b/SBOX[11].sbox/z[12] , \b/SBOX[11].sbox/z[13] ,
         \b/SBOX[11].sbox/z[14] , \b/SBOX[11].sbox/z[15] ,
         \b/SBOX[11].sbox/z[16] , \b/SBOX[11].sbox/z[17] ,
         \b/SBOX[11].sbox/t[2] , \b/SBOX[11].sbox/t[3] ,
         \b/SBOX[11].sbox/t[5] , \b/SBOX[11].sbox/t[7] ,
         \b/SBOX[11].sbox/t[8] , \b/SBOX[11].sbox/t[10] ,
         \b/SBOX[11].sbox/t[12] , \b/SBOX[11].sbox/t[13] ,
         \b/SBOX[11].sbox/t[15] , \b/SBOX[11].sbox/t[21] ,
         \b/SBOX[11].sbox/t[23] , \b/SBOX[11].sbox/t[24] ,
         \b/SBOX[11].sbox/t[25] , \b/SBOX[11].sbox/t[26] ,
         \b/SBOX[11].sbox/t[27] , \b/SBOX[11].sbox/t[28] ,
         \b/SBOX[11].sbox/t[29] , \b/SBOX[11].sbox/t[30] ,
         \b/SBOX[11].sbox/t[31] , \b/SBOX[11].sbox/t[32] ,
         \b/SBOX[11].sbox/t[33] , \b/SBOX[11].sbox/t[36] ,
         \b/SBOX[11].sbox/t[37] , \b/SBOX[11].sbox/t[38] ,
         \b/SBOX[11].sbox/t[39] , \b/SBOX[11].sbox/t[40] ,
         \b/SBOX[11].sbox/t[41] , \b/SBOX[11].sbox/t[42] ,
         \b/SBOX[11].sbox/t[43] , \b/SBOX[11].sbox/t[44] ,
         \b/SBOX[11].sbox/t[45] , \b/SBOX[11].sbox/y[1] ,
         \b/SBOX[11].sbox/y[2] , \b/SBOX[11].sbox/y[3] ,
         \b/SBOX[11].sbox/y[4] , \b/SBOX[11].sbox/y[5] ,
         \b/SBOX[11].sbox/y[6] , \b/SBOX[11].sbox/y[7] ,
         \b/SBOX[11].sbox/y[10] , \b/SBOX[11].sbox/y[11] ,
         \b/SBOX[11].sbox/y[12] , \b/SBOX[11].sbox/y[15] ,
         \b/SBOX[11].sbox/y[16] , \b/SBOX[11].sbox/y[17] ,
         \b/SBOX[10].sbox/z[0] , \b/SBOX[10].sbox/z[1] ,
         \b/SBOX[10].sbox/z[2] , \b/SBOX[10].sbox/z[3] ,
         \b/SBOX[10].sbox/z[4] , \b/SBOX[10].sbox/z[5] ,
         \b/SBOX[10].sbox/z[6] , \b/SBOX[10].sbox/z[7] ,
         \b/SBOX[10].sbox/z[8] , \b/SBOX[10].sbox/z[9] ,
         \b/SBOX[10].sbox/z[10] , \b/SBOX[10].sbox/z[11] ,
         \b/SBOX[10].sbox/z[12] , \b/SBOX[10].sbox/z[13] ,
         \b/SBOX[10].sbox/z[14] , \b/SBOX[10].sbox/z[15] ,
         \b/SBOX[10].sbox/z[16] , \b/SBOX[10].sbox/z[17] ,
         \b/SBOX[10].sbox/t[2] , \b/SBOX[10].sbox/t[3] ,
         \b/SBOX[10].sbox/t[5] , \b/SBOX[10].sbox/t[7] ,
         \b/SBOX[10].sbox/t[8] , \b/SBOX[10].sbox/t[10] ,
         \b/SBOX[10].sbox/t[12] , \b/SBOX[10].sbox/t[13] ,
         \b/SBOX[10].sbox/t[15] , \b/SBOX[10].sbox/t[21] ,
         \b/SBOX[10].sbox/t[23] , \b/SBOX[10].sbox/t[24] ,
         \b/SBOX[10].sbox/t[25] , \b/SBOX[10].sbox/t[26] ,
         \b/SBOX[10].sbox/t[27] , \b/SBOX[10].sbox/t[28] ,
         \b/SBOX[10].sbox/t[29] , \b/SBOX[10].sbox/t[30] ,
         \b/SBOX[10].sbox/t[31] , \b/SBOX[10].sbox/t[32] ,
         \b/SBOX[10].sbox/t[33] , \b/SBOX[10].sbox/t[36] ,
         \b/SBOX[10].sbox/t[37] , \b/SBOX[10].sbox/t[38] ,
         \b/SBOX[10].sbox/t[39] , \b/SBOX[10].sbox/t[40] ,
         \b/SBOX[10].sbox/t[41] , \b/SBOX[10].sbox/t[42] ,
         \b/SBOX[10].sbox/t[43] , \b/SBOX[10].sbox/t[44] ,
         \b/SBOX[10].sbox/t[45] , \b/SBOX[10].sbox/y[1] ,
         \b/SBOX[10].sbox/y[2] , \b/SBOX[10].sbox/y[3] ,
         \b/SBOX[10].sbox/y[4] , \b/SBOX[10].sbox/y[5] ,
         \b/SBOX[10].sbox/y[6] , \b/SBOX[10].sbox/y[7] ,
         \b/SBOX[10].sbox/y[10] , \b/SBOX[10].sbox/y[11] ,
         \b/SBOX[10].sbox/y[12] , \b/SBOX[10].sbox/y[15] ,
         \b/SBOX[10].sbox/y[16] , \b/SBOX[10].sbox/y[17] ,
         \b/SBOX[9].sbox/z[0] , \b/SBOX[9].sbox/z[1] , \b/SBOX[9].sbox/z[2] ,
         \b/SBOX[9].sbox/z[3] , \b/SBOX[9].sbox/z[4] , \b/SBOX[9].sbox/z[5] ,
         \b/SBOX[9].sbox/z[6] , \b/SBOX[9].sbox/z[7] , \b/SBOX[9].sbox/z[8] ,
         \b/SBOX[9].sbox/z[9] , \b/SBOX[9].sbox/z[10] , \b/SBOX[9].sbox/z[11] ,
         \b/SBOX[9].sbox/z[12] , \b/SBOX[9].sbox/z[13] ,
         \b/SBOX[9].sbox/z[14] , \b/SBOX[9].sbox/z[15] ,
         \b/SBOX[9].sbox/z[16] , \b/SBOX[9].sbox/z[17] , \b/SBOX[9].sbox/t[2] ,
         \b/SBOX[9].sbox/t[3] , \b/SBOX[9].sbox/t[5] , \b/SBOX[9].sbox/t[7] ,
         \b/SBOX[9].sbox/t[8] , \b/SBOX[9].sbox/t[10] , \b/SBOX[9].sbox/t[12] ,
         \b/SBOX[9].sbox/t[13] , \b/SBOX[9].sbox/t[15] ,
         \b/SBOX[9].sbox/t[21] , \b/SBOX[9].sbox/t[23] ,
         \b/SBOX[9].sbox/t[24] , \b/SBOX[9].sbox/t[25] ,
         \b/SBOX[9].sbox/t[26] , \b/SBOX[9].sbox/t[27] ,
         \b/SBOX[9].sbox/t[28] , \b/SBOX[9].sbox/t[29] ,
         \b/SBOX[9].sbox/t[30] , \b/SBOX[9].sbox/t[31] ,
         \b/SBOX[9].sbox/t[32] , \b/SBOX[9].sbox/t[33] ,
         \b/SBOX[9].sbox/t[36] , \b/SBOX[9].sbox/t[37] ,
         \b/SBOX[9].sbox/t[38] , \b/SBOX[9].sbox/t[39] ,
         \b/SBOX[9].sbox/t[40] , \b/SBOX[9].sbox/t[41] ,
         \b/SBOX[9].sbox/t[42] , \b/SBOX[9].sbox/t[43] ,
         \b/SBOX[9].sbox/t[44] , \b/SBOX[9].sbox/t[45] , \b/SBOX[9].sbox/y[1] ,
         \b/SBOX[9].sbox/y[2] , \b/SBOX[9].sbox/y[3] , \b/SBOX[9].sbox/y[4] ,
         \b/SBOX[9].sbox/y[5] , \b/SBOX[9].sbox/y[6] , \b/SBOX[9].sbox/y[7] ,
         \b/SBOX[9].sbox/y[10] , \b/SBOX[9].sbox/y[11] ,
         \b/SBOX[9].sbox/y[12] , \b/SBOX[9].sbox/y[15] ,
         \b/SBOX[9].sbox/y[16] , \b/SBOX[9].sbox/y[17] , \b/SBOX[8].sbox/z[0] ,
         \b/SBOX[8].sbox/z[1] , \b/SBOX[8].sbox/z[2] , \b/SBOX[8].sbox/z[3] ,
         \b/SBOX[8].sbox/z[4] , \b/SBOX[8].sbox/z[5] , \b/SBOX[8].sbox/z[6] ,
         \b/SBOX[8].sbox/z[7] , \b/SBOX[8].sbox/z[8] , \b/SBOX[8].sbox/z[9] ,
         \b/SBOX[8].sbox/z[10] , \b/SBOX[8].sbox/z[11] ,
         \b/SBOX[8].sbox/z[12] , \b/SBOX[8].sbox/z[13] ,
         \b/SBOX[8].sbox/z[14] , \b/SBOX[8].sbox/z[15] ,
         \b/SBOX[8].sbox/z[16] , \b/SBOX[8].sbox/z[17] , \b/SBOX[8].sbox/t[2] ,
         \b/SBOX[8].sbox/t[3] , \b/SBOX[8].sbox/t[5] , \b/SBOX[8].sbox/t[7] ,
         \b/SBOX[8].sbox/t[8] , \b/SBOX[8].sbox/t[10] , \b/SBOX[8].sbox/t[12] ,
         \b/SBOX[8].sbox/t[13] , \b/SBOX[8].sbox/t[15] ,
         \b/SBOX[8].sbox/t[21] , \b/SBOX[8].sbox/t[23] ,
         \b/SBOX[8].sbox/t[24] , \b/SBOX[8].sbox/t[25] ,
         \b/SBOX[8].sbox/t[26] , \b/SBOX[8].sbox/t[27] ,
         \b/SBOX[8].sbox/t[28] , \b/SBOX[8].sbox/t[29] ,
         \b/SBOX[8].sbox/t[30] , \b/SBOX[8].sbox/t[31] ,
         \b/SBOX[8].sbox/t[32] , \b/SBOX[8].sbox/t[33] ,
         \b/SBOX[8].sbox/t[36] , \b/SBOX[8].sbox/t[37] ,
         \b/SBOX[8].sbox/t[38] , \b/SBOX[8].sbox/t[39] ,
         \b/SBOX[8].sbox/t[40] , \b/SBOX[8].sbox/t[41] ,
         \b/SBOX[8].sbox/t[42] , \b/SBOX[8].sbox/t[43] ,
         \b/SBOX[8].sbox/t[44] , \b/SBOX[8].sbox/t[45] , \b/SBOX[8].sbox/y[1] ,
         \b/SBOX[8].sbox/y[2] , \b/SBOX[8].sbox/y[3] , \b/SBOX[8].sbox/y[4] ,
         \b/SBOX[8].sbox/y[5] , \b/SBOX[8].sbox/y[6] , \b/SBOX[8].sbox/y[7] ,
         \b/SBOX[8].sbox/y[10] , \b/SBOX[8].sbox/y[11] ,
         \b/SBOX[8].sbox/y[12] , \b/SBOX[8].sbox/y[15] ,
         \b/SBOX[8].sbox/y[16] , \b/SBOX[8].sbox/y[17] , \b/SBOX[7].sbox/z[0] ,
         \b/SBOX[7].sbox/z[1] , \b/SBOX[7].sbox/z[2] , \b/SBOX[7].sbox/z[3] ,
         \b/SBOX[7].sbox/z[4] , \b/SBOX[7].sbox/z[5] , \b/SBOX[7].sbox/z[6] ,
         \b/SBOX[7].sbox/z[7] , \b/SBOX[7].sbox/z[8] , \b/SBOX[7].sbox/z[9] ,
         \b/SBOX[7].sbox/z[10] , \b/SBOX[7].sbox/z[11] ,
         \b/SBOX[7].sbox/z[12] , \b/SBOX[7].sbox/z[13] ,
         \b/SBOX[7].sbox/z[14] , \b/SBOX[7].sbox/z[15] ,
         \b/SBOX[7].sbox/z[16] , \b/SBOX[7].sbox/z[17] , \b/SBOX[7].sbox/t[2] ,
         \b/SBOX[7].sbox/t[3] , \b/SBOX[7].sbox/t[5] , \b/SBOX[7].sbox/t[7] ,
         \b/SBOX[7].sbox/t[8] , \b/SBOX[7].sbox/t[10] , \b/SBOX[7].sbox/t[12] ,
         \b/SBOX[7].sbox/t[13] , \b/SBOX[7].sbox/t[15] ,
         \b/SBOX[7].sbox/t[21] , \b/SBOX[7].sbox/t[23] ,
         \b/SBOX[7].sbox/t[24] , \b/SBOX[7].sbox/t[25] ,
         \b/SBOX[7].sbox/t[26] , \b/SBOX[7].sbox/t[27] ,
         \b/SBOX[7].sbox/t[28] , \b/SBOX[7].sbox/t[29] ,
         \b/SBOX[7].sbox/t[30] , \b/SBOX[7].sbox/t[31] ,
         \b/SBOX[7].sbox/t[32] , \b/SBOX[7].sbox/t[33] ,
         \b/SBOX[7].sbox/t[36] , \b/SBOX[7].sbox/t[37] ,
         \b/SBOX[7].sbox/t[38] , \b/SBOX[7].sbox/t[39] ,
         \b/SBOX[7].sbox/t[40] , \b/SBOX[7].sbox/t[41] ,
         \b/SBOX[7].sbox/t[42] , \b/SBOX[7].sbox/t[43] ,
         \b/SBOX[7].sbox/t[44] , \b/SBOX[7].sbox/t[45] , \b/SBOX[7].sbox/y[1] ,
         \b/SBOX[7].sbox/y[2] , \b/SBOX[7].sbox/y[3] , \b/SBOX[7].sbox/y[4] ,
         \b/SBOX[7].sbox/y[5] , \b/SBOX[7].sbox/y[6] , \b/SBOX[7].sbox/y[7] ,
         \b/SBOX[7].sbox/y[10] , \b/SBOX[7].sbox/y[11] ,
         \b/SBOX[7].sbox/y[12] , \b/SBOX[7].sbox/y[15] ,
         \b/SBOX[7].sbox/y[16] , \b/SBOX[7].sbox/y[17] , \b/SBOX[6].sbox/z[0] ,
         \b/SBOX[6].sbox/z[1] , \b/SBOX[6].sbox/z[2] , \b/SBOX[6].sbox/z[3] ,
         \b/SBOX[6].sbox/z[4] , \b/SBOX[6].sbox/z[5] , \b/SBOX[6].sbox/z[6] ,
         \b/SBOX[6].sbox/z[7] , \b/SBOX[6].sbox/z[8] , \b/SBOX[6].sbox/z[9] ,
         \b/SBOX[6].sbox/z[10] , \b/SBOX[6].sbox/z[11] ,
         \b/SBOX[6].sbox/z[12] , \b/SBOX[6].sbox/z[13] ,
         \b/SBOX[6].sbox/z[14] , \b/SBOX[6].sbox/z[15] ,
         \b/SBOX[6].sbox/z[16] , \b/SBOX[6].sbox/z[17] , \b/SBOX[6].sbox/t[2] ,
         \b/SBOX[6].sbox/t[3] , \b/SBOX[6].sbox/t[5] , \b/SBOX[6].sbox/t[7] ,
         \b/SBOX[6].sbox/t[8] , \b/SBOX[6].sbox/t[10] , \b/SBOX[6].sbox/t[12] ,
         \b/SBOX[6].sbox/t[13] , \b/SBOX[6].sbox/t[15] ,
         \b/SBOX[6].sbox/t[21] , \b/SBOX[6].sbox/t[23] ,
         \b/SBOX[6].sbox/t[24] , \b/SBOX[6].sbox/t[25] ,
         \b/SBOX[6].sbox/t[26] , \b/SBOX[6].sbox/t[27] ,
         \b/SBOX[6].sbox/t[28] , \b/SBOX[6].sbox/t[29] ,
         \b/SBOX[6].sbox/t[30] , \b/SBOX[6].sbox/t[31] ,
         \b/SBOX[6].sbox/t[32] , \b/SBOX[6].sbox/t[33] ,
         \b/SBOX[6].sbox/t[36] , \b/SBOX[6].sbox/t[37] ,
         \b/SBOX[6].sbox/t[38] , \b/SBOX[6].sbox/t[39] ,
         \b/SBOX[6].sbox/t[40] , \b/SBOX[6].sbox/t[41] ,
         \b/SBOX[6].sbox/t[42] , \b/SBOX[6].sbox/t[43] ,
         \b/SBOX[6].sbox/t[44] , \b/SBOX[6].sbox/t[45] , \b/SBOX[6].sbox/y[1] ,
         \b/SBOX[6].sbox/y[2] , \b/SBOX[6].sbox/y[3] , \b/SBOX[6].sbox/y[4] ,
         \b/SBOX[6].sbox/y[5] , \b/SBOX[6].sbox/y[6] , \b/SBOX[6].sbox/y[7] ,
         \b/SBOX[6].sbox/y[10] , \b/SBOX[6].sbox/y[11] ,
         \b/SBOX[6].sbox/y[12] , \b/SBOX[6].sbox/y[15] ,
         \b/SBOX[6].sbox/y[16] , \b/SBOX[6].sbox/y[17] , \b/SBOX[5].sbox/z[0] ,
         \b/SBOX[5].sbox/z[1] , \b/SBOX[5].sbox/z[2] , \b/SBOX[5].sbox/z[3] ,
         \b/SBOX[5].sbox/z[4] , \b/SBOX[5].sbox/z[5] , \b/SBOX[5].sbox/z[6] ,
         \b/SBOX[5].sbox/z[7] , \b/SBOX[5].sbox/z[8] , \b/SBOX[5].sbox/z[9] ,
         \b/SBOX[5].sbox/z[10] , \b/SBOX[5].sbox/z[11] ,
         \b/SBOX[5].sbox/z[12] , \b/SBOX[5].sbox/z[13] ,
         \b/SBOX[5].sbox/z[14] , \b/SBOX[5].sbox/z[15] ,
         \b/SBOX[5].sbox/z[16] , \b/SBOX[5].sbox/z[17] , \b/SBOX[5].sbox/t[2] ,
         \b/SBOX[5].sbox/t[3] , \b/SBOX[5].sbox/t[5] , \b/SBOX[5].sbox/t[7] ,
         \b/SBOX[5].sbox/t[8] , \b/SBOX[5].sbox/t[10] , \b/SBOX[5].sbox/t[12] ,
         \b/SBOX[5].sbox/t[13] , \b/SBOX[5].sbox/t[15] ,
         \b/SBOX[5].sbox/t[21] , \b/SBOX[5].sbox/t[23] ,
         \b/SBOX[5].sbox/t[24] , \b/SBOX[5].sbox/t[25] ,
         \b/SBOX[5].sbox/t[26] , \b/SBOX[5].sbox/t[27] ,
         \b/SBOX[5].sbox/t[28] , \b/SBOX[5].sbox/t[29] ,
         \b/SBOX[5].sbox/t[30] , \b/SBOX[5].sbox/t[31] ,
         \b/SBOX[5].sbox/t[32] , \b/SBOX[5].sbox/t[33] ,
         \b/SBOX[5].sbox/t[36] , \b/SBOX[5].sbox/t[37] ,
         \b/SBOX[5].sbox/t[38] , \b/SBOX[5].sbox/t[39] ,
         \b/SBOX[5].sbox/t[40] , \b/SBOX[5].sbox/t[41] ,
         \b/SBOX[5].sbox/t[42] , \b/SBOX[5].sbox/t[43] ,
         \b/SBOX[5].sbox/t[44] , \b/SBOX[5].sbox/t[45] , \b/SBOX[5].sbox/y[1] ,
         \b/SBOX[5].sbox/y[2] , \b/SBOX[5].sbox/y[3] , \b/SBOX[5].sbox/y[4] ,
         \b/SBOX[5].sbox/y[5] , \b/SBOX[5].sbox/y[6] , \b/SBOX[5].sbox/y[7] ,
         \b/SBOX[5].sbox/y[10] , \b/SBOX[5].sbox/y[11] ,
         \b/SBOX[5].sbox/y[12] , \b/SBOX[5].sbox/y[15] ,
         \b/SBOX[5].sbox/y[16] , \b/SBOX[5].sbox/y[17] , \b/SBOX[4].sbox/z[0] ,
         \b/SBOX[4].sbox/z[1] , \b/SBOX[4].sbox/z[2] , \b/SBOX[4].sbox/z[3] ,
         \b/SBOX[4].sbox/z[4] , \b/SBOX[4].sbox/z[5] , \b/SBOX[4].sbox/z[6] ,
         \b/SBOX[4].sbox/z[7] , \b/SBOX[4].sbox/z[8] , \b/SBOX[4].sbox/z[9] ,
         \b/SBOX[4].sbox/z[10] , \b/SBOX[4].sbox/z[11] ,
         \b/SBOX[4].sbox/z[12] , \b/SBOX[4].sbox/z[13] ,
         \b/SBOX[4].sbox/z[14] , \b/SBOX[4].sbox/z[15] ,
         \b/SBOX[4].sbox/z[16] , \b/SBOX[4].sbox/z[17] , \b/SBOX[4].sbox/t[2] ,
         \b/SBOX[4].sbox/t[3] , \b/SBOX[4].sbox/t[5] , \b/SBOX[4].sbox/t[7] ,
         \b/SBOX[4].sbox/t[8] , \b/SBOX[4].sbox/t[10] , \b/SBOX[4].sbox/t[12] ,
         \b/SBOX[4].sbox/t[13] , \b/SBOX[4].sbox/t[15] ,
         \b/SBOX[4].sbox/t[21] , \b/SBOX[4].sbox/t[23] ,
         \b/SBOX[4].sbox/t[24] , \b/SBOX[4].sbox/t[25] ,
         \b/SBOX[4].sbox/t[26] , \b/SBOX[4].sbox/t[27] ,
         \b/SBOX[4].sbox/t[28] , \b/SBOX[4].sbox/t[29] ,
         \b/SBOX[4].sbox/t[30] , \b/SBOX[4].sbox/t[31] ,
         \b/SBOX[4].sbox/t[32] , \b/SBOX[4].sbox/t[33] ,
         \b/SBOX[4].sbox/t[36] , \b/SBOX[4].sbox/t[37] ,
         \b/SBOX[4].sbox/t[38] , \b/SBOX[4].sbox/t[39] ,
         \b/SBOX[4].sbox/t[40] , \b/SBOX[4].sbox/t[41] ,
         \b/SBOX[4].sbox/t[42] , \b/SBOX[4].sbox/t[43] ,
         \b/SBOX[4].sbox/t[44] , \b/SBOX[4].sbox/t[45] , \b/SBOX[4].sbox/y[1] ,
         \b/SBOX[4].sbox/y[2] , \b/SBOX[4].sbox/y[3] , \b/SBOX[4].sbox/y[4] ,
         \b/SBOX[4].sbox/y[5] , \b/SBOX[4].sbox/y[6] , \b/SBOX[4].sbox/y[7] ,
         \b/SBOX[4].sbox/y[10] , \b/SBOX[4].sbox/y[11] ,
         \b/SBOX[4].sbox/y[12] , \b/SBOX[4].sbox/y[15] ,
         \b/SBOX[4].sbox/y[16] , \b/SBOX[4].sbox/y[17] , \b/SBOX[3].sbox/z[0] ,
         \b/SBOX[3].sbox/z[1] , \b/SBOX[3].sbox/z[2] , \b/SBOX[3].sbox/z[3] ,
         \b/SBOX[3].sbox/z[4] , \b/SBOX[3].sbox/z[5] , \b/SBOX[3].sbox/z[6] ,
         \b/SBOX[3].sbox/z[7] , \b/SBOX[3].sbox/z[8] , \b/SBOX[3].sbox/z[9] ,
         \b/SBOX[3].sbox/z[10] , \b/SBOX[3].sbox/z[11] ,
         \b/SBOX[3].sbox/z[12] , \b/SBOX[3].sbox/z[13] ,
         \b/SBOX[3].sbox/z[14] , \b/SBOX[3].sbox/z[15] ,
         \b/SBOX[3].sbox/z[16] , \b/SBOX[3].sbox/z[17] , \b/SBOX[3].sbox/t[2] ,
         \b/SBOX[3].sbox/t[3] , \b/SBOX[3].sbox/t[5] , \b/SBOX[3].sbox/t[7] ,
         \b/SBOX[3].sbox/t[8] , \b/SBOX[3].sbox/t[10] , \b/SBOX[3].sbox/t[12] ,
         \b/SBOX[3].sbox/t[13] , \b/SBOX[3].sbox/t[15] ,
         \b/SBOX[3].sbox/t[21] , \b/SBOX[3].sbox/t[23] ,
         \b/SBOX[3].sbox/t[24] , \b/SBOX[3].sbox/t[25] ,
         \b/SBOX[3].sbox/t[26] , \b/SBOX[3].sbox/t[27] ,
         \b/SBOX[3].sbox/t[28] , \b/SBOX[3].sbox/t[29] ,
         \b/SBOX[3].sbox/t[30] , \b/SBOX[3].sbox/t[31] ,
         \b/SBOX[3].sbox/t[32] , \b/SBOX[3].sbox/t[33] ,
         \b/SBOX[3].sbox/t[36] , \b/SBOX[3].sbox/t[37] ,
         \b/SBOX[3].sbox/t[38] , \b/SBOX[3].sbox/t[39] ,
         \b/SBOX[3].sbox/t[40] , \b/SBOX[3].sbox/t[41] ,
         \b/SBOX[3].sbox/t[42] , \b/SBOX[3].sbox/t[43] ,
         \b/SBOX[3].sbox/t[44] , \b/SBOX[3].sbox/t[45] , \b/SBOX[3].sbox/y[1] ,
         \b/SBOX[3].sbox/y[2] , \b/SBOX[3].sbox/y[3] , \b/SBOX[3].sbox/y[4] ,
         \b/SBOX[3].sbox/y[5] , \b/SBOX[3].sbox/y[6] , \b/SBOX[3].sbox/y[7] ,
         \b/SBOX[3].sbox/y[10] , \b/SBOX[3].sbox/y[11] ,
         \b/SBOX[3].sbox/y[12] , \b/SBOX[3].sbox/y[15] ,
         \b/SBOX[3].sbox/y[16] , \b/SBOX[3].sbox/y[17] , \b/SBOX[2].sbox/z[0] ,
         \b/SBOX[2].sbox/z[1] , \b/SBOX[2].sbox/z[2] , \b/SBOX[2].sbox/z[3] ,
         \b/SBOX[2].sbox/z[4] , \b/SBOX[2].sbox/z[5] , \b/SBOX[2].sbox/z[6] ,
         \b/SBOX[2].sbox/z[7] , \b/SBOX[2].sbox/z[8] , \b/SBOX[2].sbox/z[9] ,
         \b/SBOX[2].sbox/z[10] , \b/SBOX[2].sbox/z[11] ,
         \b/SBOX[2].sbox/z[12] , \b/SBOX[2].sbox/z[13] ,
         \b/SBOX[2].sbox/z[14] , \b/SBOX[2].sbox/z[15] ,
         \b/SBOX[2].sbox/z[16] , \b/SBOX[2].sbox/z[17] , \b/SBOX[2].sbox/t[2] ,
         \b/SBOX[2].sbox/t[3] , \b/SBOX[2].sbox/t[5] , \b/SBOX[2].sbox/t[7] ,
         \b/SBOX[2].sbox/t[8] , \b/SBOX[2].sbox/t[10] , \b/SBOX[2].sbox/t[12] ,
         \b/SBOX[2].sbox/t[13] , \b/SBOX[2].sbox/t[15] ,
         \b/SBOX[2].sbox/t[21] , \b/SBOX[2].sbox/t[23] ,
         \b/SBOX[2].sbox/t[24] , \b/SBOX[2].sbox/t[25] ,
         \b/SBOX[2].sbox/t[26] , \b/SBOX[2].sbox/t[27] ,
         \b/SBOX[2].sbox/t[28] , \b/SBOX[2].sbox/t[29] ,
         \b/SBOX[2].sbox/t[30] , \b/SBOX[2].sbox/t[31] ,
         \b/SBOX[2].sbox/t[32] , \b/SBOX[2].sbox/t[33] ,
         \b/SBOX[2].sbox/t[36] , \b/SBOX[2].sbox/t[37] ,
         \b/SBOX[2].sbox/t[38] , \b/SBOX[2].sbox/t[39] ,
         \b/SBOX[2].sbox/t[40] , \b/SBOX[2].sbox/t[41] ,
         \b/SBOX[2].sbox/t[42] , \b/SBOX[2].sbox/t[43] ,
         \b/SBOX[2].sbox/t[44] , \b/SBOX[2].sbox/t[45] , \b/SBOX[2].sbox/y[1] ,
         \b/SBOX[2].sbox/y[2] , \b/SBOX[2].sbox/y[3] , \b/SBOX[2].sbox/y[4] ,
         \b/SBOX[2].sbox/y[5] , \b/SBOX[2].sbox/y[6] , \b/SBOX[2].sbox/y[7] ,
         \b/SBOX[2].sbox/y[10] , \b/SBOX[2].sbox/y[11] ,
         \b/SBOX[2].sbox/y[12] , \b/SBOX[2].sbox/y[15] ,
         \b/SBOX[2].sbox/y[16] , \b/SBOX[2].sbox/y[17] , \b/SBOX[1].sbox/z[0] ,
         \b/SBOX[1].sbox/z[1] , \b/SBOX[1].sbox/z[2] , \b/SBOX[1].sbox/z[3] ,
         \b/SBOX[1].sbox/z[4] , \b/SBOX[1].sbox/z[5] , \b/SBOX[1].sbox/z[6] ,
         \b/SBOX[1].sbox/z[7] , \b/SBOX[1].sbox/z[8] , \b/SBOX[1].sbox/z[9] ,
         \b/SBOX[1].sbox/z[10] , \b/SBOX[1].sbox/z[11] ,
         \b/SBOX[1].sbox/z[12] , \b/SBOX[1].sbox/z[13] ,
         \b/SBOX[1].sbox/z[14] , \b/SBOX[1].sbox/z[15] ,
         \b/SBOX[1].sbox/z[16] , \b/SBOX[1].sbox/z[17] , \b/SBOX[1].sbox/t[2] ,
         \b/SBOX[1].sbox/t[3] , \b/SBOX[1].sbox/t[5] , \b/SBOX[1].sbox/t[7] ,
         \b/SBOX[1].sbox/t[8] , \b/SBOX[1].sbox/t[10] , \b/SBOX[1].sbox/t[12] ,
         \b/SBOX[1].sbox/t[13] , \b/SBOX[1].sbox/t[15] ,
         \b/SBOX[1].sbox/t[21] , \b/SBOX[1].sbox/t[23] ,
         \b/SBOX[1].sbox/t[24] , \b/SBOX[1].sbox/t[25] ,
         \b/SBOX[1].sbox/t[26] , \b/SBOX[1].sbox/t[27] ,
         \b/SBOX[1].sbox/t[28] , \b/SBOX[1].sbox/t[29] ,
         \b/SBOX[1].sbox/t[30] , \b/SBOX[1].sbox/t[31] ,
         \b/SBOX[1].sbox/t[32] , \b/SBOX[1].sbox/t[33] ,
         \b/SBOX[1].sbox/t[36] , \b/SBOX[1].sbox/t[37] ,
         \b/SBOX[1].sbox/t[38] , \b/SBOX[1].sbox/t[39] ,
         \b/SBOX[1].sbox/t[40] , \b/SBOX[1].sbox/t[41] ,
         \b/SBOX[1].sbox/t[42] , \b/SBOX[1].sbox/t[43] ,
         \b/SBOX[1].sbox/t[44] , \b/SBOX[1].sbox/t[45] , \b/SBOX[1].sbox/y[1] ,
         \b/SBOX[1].sbox/y[2] , \b/SBOX[1].sbox/y[3] , \b/SBOX[1].sbox/y[4] ,
         \b/SBOX[1].sbox/y[5] , \b/SBOX[1].sbox/y[6] , \b/SBOX[1].sbox/y[7] ,
         \b/SBOX[1].sbox/y[10] , \b/SBOX[1].sbox/y[11] ,
         \b/SBOX[1].sbox/y[12] , \b/SBOX[1].sbox/y[15] ,
         \b/SBOX[1].sbox/y[16] , \b/SBOX[1].sbox/y[17] , n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328;
  wire   [127:0] key;
  wire   [3:0] counter;
  wire   [127:0] nextKey;
  wire   [127:0] msg;
  wire   [127:0] shift_row_out;

  DFF \counter_reg[0]  ( .D(n7), .CLK(clk), .RST(rst), .I(1'b0), .Q(counter[0]) );
  DFF \counter_reg[1]  ( .D(N5), .CLK(clk), .RST(rst), .I(1'b0), .Q(counter[1]) );
  DFF \counter_reg[2]  ( .D(N6), .CLK(clk), .RST(rst), .I(1'b0), .Q(counter[2]) );
  DFF \counter_reg[3]  ( .D(N7), .CLK(clk), .RST(rst), .I(1'b0), .Q(counter[3]) );
  DFF \key_reg[0]  ( .D(nextKey[0]), .CLK(clk), .RST(rst), .I(g_init[0]), .Q(
        key[0]) );
  DFF \key_reg[1]  ( .D(nextKey[1]), .CLK(clk), .RST(rst), .I(g_init[1]), .Q(
        key[1]) );
  DFF \key_reg[2]  ( .D(nextKey[2]), .CLK(clk), .RST(rst), .I(g_init[2]), .Q(
        key[2]) );
  DFF \key_reg[3]  ( .D(nextKey[3]), .CLK(clk), .RST(rst), .I(g_init[3]), .Q(
        key[3]) );
  DFF \key_reg[4]  ( .D(nextKey[4]), .CLK(clk), .RST(rst), .I(g_init[4]), .Q(
        key[4]) );
  DFF \key_reg[5]  ( .D(nextKey[5]), .CLK(clk), .RST(rst), .I(g_init[5]), .Q(
        key[5]) );
  DFF \key_reg[6]  ( .D(nextKey[6]), .CLK(clk), .RST(rst), .I(g_init[6]), .Q(
        key[6]) );
  DFF \key_reg[7]  ( .D(nextKey[7]), .CLK(clk), .RST(rst), .I(g_init[7]), .Q(
        key[7]) );
  DFF \key_reg[8]  ( .D(nextKey[8]), .CLK(clk), .RST(rst), .I(g_init[8]), .Q(
        key[8]) );
  DFF \key_reg[9]  ( .D(nextKey[9]), .CLK(clk), .RST(rst), .I(g_init[9]), .Q(
        key[9]) );
  DFF \key_reg[10]  ( .D(nextKey[10]), .CLK(clk), .RST(rst), .I(g_init[10]), 
        .Q(key[10]) );
  DFF \key_reg[11]  ( .D(nextKey[11]), .CLK(clk), .RST(rst), .I(g_init[11]), 
        .Q(key[11]) );
  DFF \key_reg[12]  ( .D(nextKey[12]), .CLK(clk), .RST(rst), .I(g_init[12]), 
        .Q(key[12]) );
  DFF \key_reg[13]  ( .D(nextKey[13]), .CLK(clk), .RST(rst), .I(g_init[13]), 
        .Q(key[13]) );
  DFF \key_reg[14]  ( .D(nextKey[14]), .CLK(clk), .RST(rst), .I(g_init[14]), 
        .Q(key[14]) );
  DFF \key_reg[15]  ( .D(nextKey[15]), .CLK(clk), .RST(rst), .I(g_init[15]), 
        .Q(key[15]) );
  DFF \key_reg[16]  ( .D(nextKey[16]), .CLK(clk), .RST(rst), .I(g_init[16]), 
        .Q(key[16]) );
  DFF \key_reg[17]  ( .D(nextKey[17]), .CLK(clk), .RST(rst), .I(g_init[17]), 
        .Q(key[17]) );
  DFF \key_reg[18]  ( .D(nextKey[18]), .CLK(clk), .RST(rst), .I(g_init[18]), 
        .Q(key[18]) );
  DFF \key_reg[19]  ( .D(nextKey[19]), .CLK(clk), .RST(rst), .I(g_init[19]), 
        .Q(key[19]) );
  DFF \key_reg[20]  ( .D(nextKey[20]), .CLK(clk), .RST(rst), .I(g_init[20]), 
        .Q(key[20]) );
  DFF \key_reg[21]  ( .D(nextKey[21]), .CLK(clk), .RST(rst), .I(g_init[21]), 
        .Q(key[21]) );
  DFF \key_reg[22]  ( .D(nextKey[22]), .CLK(clk), .RST(rst), .I(g_init[22]), 
        .Q(key[22]) );
  DFF \key_reg[23]  ( .D(nextKey[23]), .CLK(clk), .RST(rst), .I(g_init[23]), 
        .Q(key[23]) );
  DFF \key_reg[24]  ( .D(nextKey[24]), .CLK(clk), .RST(rst), .I(g_init[24]), 
        .Q(key[24]) );
  DFF \key_reg[25]  ( .D(nextKey[25]), .CLK(clk), .RST(rst), .I(g_init[25]), 
        .Q(key[25]) );
  DFF \key_reg[26]  ( .D(nextKey[26]), .CLK(clk), .RST(rst), .I(g_init[26]), 
        .Q(key[26]) );
  DFF \key_reg[27]  ( .D(nextKey[27]), .CLK(clk), .RST(rst), .I(g_init[27]), 
        .Q(key[27]) );
  DFF \key_reg[28]  ( .D(nextKey[28]), .CLK(clk), .RST(rst), .I(g_init[28]), 
        .Q(key[28]) );
  DFF \key_reg[29]  ( .D(nextKey[29]), .CLK(clk), .RST(rst), .I(g_init[29]), 
        .Q(key[29]) );
  DFF \key_reg[30]  ( .D(nextKey[30]), .CLK(clk), .RST(rst), .I(g_init[30]), 
        .Q(key[30]) );
  DFF \key_reg[31]  ( .D(nextKey[31]), .CLK(clk), .RST(rst), .I(g_init[31]), 
        .Q(key[31]) );
  DFF \key_reg[32]  ( .D(nextKey[32]), .CLK(clk), .RST(rst), .I(g_init[32]), 
        .Q(key[32]) );
  DFF \key_reg[33]  ( .D(nextKey[33]), .CLK(clk), .RST(rst), .I(g_init[33]), 
        .Q(key[33]) );
  DFF \key_reg[34]  ( .D(nextKey[34]), .CLK(clk), .RST(rst), .I(g_init[34]), 
        .Q(key[34]) );
  DFF \key_reg[35]  ( .D(nextKey[35]), .CLK(clk), .RST(rst), .I(g_init[35]), 
        .Q(key[35]) );
  DFF \key_reg[36]  ( .D(nextKey[36]), .CLK(clk), .RST(rst), .I(g_init[36]), 
        .Q(key[36]) );
  DFF \key_reg[37]  ( .D(nextKey[37]), .CLK(clk), .RST(rst), .I(g_init[37]), 
        .Q(key[37]) );
  DFF \key_reg[38]  ( .D(nextKey[38]), .CLK(clk), .RST(rst), .I(g_init[38]), 
        .Q(key[38]) );
  DFF \key_reg[39]  ( .D(nextKey[39]), .CLK(clk), .RST(rst), .I(g_init[39]), 
        .Q(key[39]) );
  DFF \key_reg[40]  ( .D(nextKey[40]), .CLK(clk), .RST(rst), .I(g_init[40]), 
        .Q(key[40]) );
  DFF \key_reg[41]  ( .D(nextKey[41]), .CLK(clk), .RST(rst), .I(g_init[41]), 
        .Q(key[41]) );
  DFF \key_reg[42]  ( .D(nextKey[42]), .CLK(clk), .RST(rst), .I(g_init[42]), 
        .Q(key[42]) );
  DFF \key_reg[43]  ( .D(nextKey[43]), .CLK(clk), .RST(rst), .I(g_init[43]), 
        .Q(key[43]) );
  DFF \key_reg[44]  ( .D(nextKey[44]), .CLK(clk), .RST(rst), .I(g_init[44]), 
        .Q(key[44]) );
  DFF \key_reg[45]  ( .D(nextKey[45]), .CLK(clk), .RST(rst), .I(g_init[45]), 
        .Q(key[45]) );
  DFF \key_reg[46]  ( .D(nextKey[46]), .CLK(clk), .RST(rst), .I(g_init[46]), 
        .Q(key[46]) );
  DFF \key_reg[47]  ( .D(nextKey[47]), .CLK(clk), .RST(rst), .I(g_init[47]), 
        .Q(key[47]) );
  DFF \key_reg[48]  ( .D(nextKey[48]), .CLK(clk), .RST(rst), .I(g_init[48]), 
        .Q(key[48]) );
  DFF \key_reg[49]  ( .D(nextKey[49]), .CLK(clk), .RST(rst), .I(g_init[49]), 
        .Q(key[49]) );
  DFF \key_reg[50]  ( .D(nextKey[50]), .CLK(clk), .RST(rst), .I(g_init[50]), 
        .Q(key[50]) );
  DFF \key_reg[51]  ( .D(nextKey[51]), .CLK(clk), .RST(rst), .I(g_init[51]), 
        .Q(key[51]) );
  DFF \key_reg[52]  ( .D(nextKey[52]), .CLK(clk), .RST(rst), .I(g_init[52]), 
        .Q(key[52]) );
  DFF \key_reg[53]  ( .D(nextKey[53]), .CLK(clk), .RST(rst), .I(g_init[53]), 
        .Q(key[53]) );
  DFF \key_reg[54]  ( .D(nextKey[54]), .CLK(clk), .RST(rst), .I(g_init[54]), 
        .Q(key[54]) );
  DFF \key_reg[55]  ( .D(nextKey[55]), .CLK(clk), .RST(rst), .I(g_init[55]), 
        .Q(key[55]) );
  DFF \key_reg[56]  ( .D(nextKey[56]), .CLK(clk), .RST(rst), .I(g_init[56]), 
        .Q(key[56]) );
  DFF \key_reg[57]  ( .D(nextKey[57]), .CLK(clk), .RST(rst), .I(g_init[57]), 
        .Q(key[57]) );
  DFF \key_reg[58]  ( .D(nextKey[58]), .CLK(clk), .RST(rst), .I(g_init[58]), 
        .Q(key[58]) );
  DFF \key_reg[59]  ( .D(nextKey[59]), .CLK(clk), .RST(rst), .I(g_init[59]), 
        .Q(key[59]) );
  DFF \key_reg[60]  ( .D(nextKey[60]), .CLK(clk), .RST(rst), .I(g_init[60]), 
        .Q(key[60]) );
  DFF \key_reg[61]  ( .D(nextKey[61]), .CLK(clk), .RST(rst), .I(g_init[61]), 
        .Q(key[61]) );
  DFF \key_reg[62]  ( .D(nextKey[62]), .CLK(clk), .RST(rst), .I(g_init[62]), 
        .Q(key[62]) );
  DFF \key_reg[63]  ( .D(nextKey[63]), .CLK(clk), .RST(rst), .I(g_init[63]), 
        .Q(key[63]) );
  DFF \key_reg[64]  ( .D(nextKey[64]), .CLK(clk), .RST(rst), .I(g_init[64]), 
        .Q(key[64]) );
  DFF \key_reg[65]  ( .D(nextKey[65]), .CLK(clk), .RST(rst), .I(g_init[65]), 
        .Q(key[65]) );
  DFF \key_reg[66]  ( .D(nextKey[66]), .CLK(clk), .RST(rst), .I(g_init[66]), 
        .Q(key[66]) );
  DFF \key_reg[67]  ( .D(nextKey[67]), .CLK(clk), .RST(rst), .I(g_init[67]), 
        .Q(key[67]) );
  DFF \key_reg[68]  ( .D(nextKey[68]), .CLK(clk), .RST(rst), .I(g_init[68]), 
        .Q(key[68]) );
  DFF \key_reg[69]  ( .D(nextKey[69]), .CLK(clk), .RST(rst), .I(g_init[69]), 
        .Q(key[69]) );
  DFF \key_reg[70]  ( .D(nextKey[70]), .CLK(clk), .RST(rst), .I(g_init[70]), 
        .Q(key[70]) );
  DFF \key_reg[71]  ( .D(nextKey[71]), .CLK(clk), .RST(rst), .I(g_init[71]), 
        .Q(key[71]) );
  DFF \key_reg[72]  ( .D(nextKey[72]), .CLK(clk), .RST(rst), .I(g_init[72]), 
        .Q(key[72]) );
  DFF \key_reg[73]  ( .D(nextKey[73]), .CLK(clk), .RST(rst), .I(g_init[73]), 
        .Q(key[73]) );
  DFF \key_reg[74]  ( .D(nextKey[74]), .CLK(clk), .RST(rst), .I(g_init[74]), 
        .Q(key[74]) );
  DFF \key_reg[75]  ( .D(nextKey[75]), .CLK(clk), .RST(rst), .I(g_init[75]), 
        .Q(key[75]) );
  DFF \key_reg[76]  ( .D(nextKey[76]), .CLK(clk), .RST(rst), .I(g_init[76]), 
        .Q(key[76]) );
  DFF \key_reg[77]  ( .D(nextKey[77]), .CLK(clk), .RST(rst), .I(g_init[77]), 
        .Q(key[77]) );
  DFF \key_reg[78]  ( .D(nextKey[78]), .CLK(clk), .RST(rst), .I(g_init[78]), 
        .Q(key[78]) );
  DFF \key_reg[79]  ( .D(nextKey[79]), .CLK(clk), .RST(rst), .I(g_init[79]), 
        .Q(key[79]) );
  DFF \key_reg[80]  ( .D(nextKey[80]), .CLK(clk), .RST(rst), .I(g_init[80]), 
        .Q(key[80]) );
  DFF \key_reg[81]  ( .D(nextKey[81]), .CLK(clk), .RST(rst), .I(g_init[81]), 
        .Q(key[81]) );
  DFF \key_reg[82]  ( .D(nextKey[82]), .CLK(clk), .RST(rst), .I(g_init[82]), 
        .Q(key[82]) );
  DFF \key_reg[83]  ( .D(nextKey[83]), .CLK(clk), .RST(rst), .I(g_init[83]), 
        .Q(key[83]) );
  DFF \key_reg[84]  ( .D(nextKey[84]), .CLK(clk), .RST(rst), .I(g_init[84]), 
        .Q(key[84]) );
  DFF \key_reg[85]  ( .D(nextKey[85]), .CLK(clk), .RST(rst), .I(g_init[85]), 
        .Q(key[85]) );
  DFF \key_reg[86]  ( .D(nextKey[86]), .CLK(clk), .RST(rst), .I(g_init[86]), 
        .Q(key[86]) );
  DFF \key_reg[87]  ( .D(nextKey[87]), .CLK(clk), .RST(rst), .I(g_init[87]), 
        .Q(key[87]) );
  DFF \key_reg[88]  ( .D(nextKey[88]), .CLK(clk), .RST(rst), .I(g_init[88]), 
        .Q(key[88]) );
  DFF \key_reg[89]  ( .D(nextKey[89]), .CLK(clk), .RST(rst), .I(g_init[89]), 
        .Q(key[89]) );
  DFF \key_reg[90]  ( .D(nextKey[90]), .CLK(clk), .RST(rst), .I(g_init[90]), 
        .Q(key[90]) );
  DFF \key_reg[91]  ( .D(nextKey[91]), .CLK(clk), .RST(rst), .I(g_init[91]), 
        .Q(key[91]) );
  DFF \key_reg[92]  ( .D(nextKey[92]), .CLK(clk), .RST(rst), .I(g_init[92]), 
        .Q(key[92]) );
  DFF \key_reg[93]  ( .D(nextKey[93]), .CLK(clk), .RST(rst), .I(g_init[93]), 
        .Q(key[93]) );
  DFF \key_reg[94]  ( .D(nextKey[94]), .CLK(clk), .RST(rst), .I(g_init[94]), 
        .Q(key[94]) );
  DFF \key_reg[95]  ( .D(nextKey[95]), .CLK(clk), .RST(rst), .I(g_init[95]), 
        .Q(key[95]) );
  DFF \key_reg[96]  ( .D(n552), .CLK(clk), .RST(rst), .I(g_init[96]), .Q(
        key[96]) );
  DFF \key_reg[97]  ( .D(n551), .CLK(clk), .RST(rst), .I(g_init[97]), .Q(
        key[97]) );
  DFF \key_reg[98]  ( .D(n550), .CLK(clk), .RST(rst), .I(g_init[98]), .Q(
        key[98]) );
  DFF \key_reg[99]  ( .D(n549), .CLK(clk), .RST(rst), .I(g_init[99]), .Q(
        key[99]) );
  DFF \key_reg[100]  ( .D(n548), .CLK(clk), .RST(rst), .I(g_init[100]), .Q(
        key[100]) );
  DFF \key_reg[101]  ( .D(n547), .CLK(clk), .RST(rst), .I(g_init[101]), .Q(
        key[101]) );
  DFF \key_reg[102]  ( .D(n546), .CLK(clk), .RST(rst), .I(g_init[102]), .Q(
        key[102]) );
  DFF \key_reg[103]  ( .D(n545), .CLK(clk), .RST(rst), .I(g_init[103]), .Q(
        key[103]) );
  DFF \key_reg[104]  ( .D(nextKey[104]), .CLK(clk), .RST(rst), .I(g_init[104]), 
        .Q(key[104]) );
  DFF \key_reg[105]  ( .D(nextKey[105]), .CLK(clk), .RST(rst), .I(g_init[105]), 
        .Q(key[105]) );
  DFF \key_reg[106]  ( .D(nextKey[106]), .CLK(clk), .RST(rst), .I(g_init[106]), 
        .Q(key[106]) );
  DFF \key_reg[107]  ( .D(nextKey[107]), .CLK(clk), .RST(rst), .I(g_init[107]), 
        .Q(key[107]) );
  DFF \key_reg[108]  ( .D(nextKey[108]), .CLK(clk), .RST(rst), .I(g_init[108]), 
        .Q(key[108]) );
  DFF \key_reg[109]  ( .D(nextKey[109]), .CLK(clk), .RST(rst), .I(g_init[109]), 
        .Q(key[109]) );
  DFF \key_reg[110]  ( .D(nextKey[110]), .CLK(clk), .RST(rst), .I(g_init[110]), 
        .Q(key[110]) );
  DFF \key_reg[111]  ( .D(nextKey[111]), .CLK(clk), .RST(rst), .I(g_init[111]), 
        .Q(key[111]) );
  DFF \key_reg[112]  ( .D(nextKey[112]), .CLK(clk), .RST(rst), .I(g_init[112]), 
        .Q(key[112]) );
  DFF \key_reg[113]  ( .D(nextKey[113]), .CLK(clk), .RST(rst), .I(g_init[113]), 
        .Q(key[113]) );
  DFF \key_reg[114]  ( .D(nextKey[114]), .CLK(clk), .RST(rst), .I(g_init[114]), 
        .Q(key[114]) );
  DFF \key_reg[115]  ( .D(nextKey[115]), .CLK(clk), .RST(rst), .I(g_init[115]), 
        .Q(key[115]) );
  DFF \key_reg[116]  ( .D(nextKey[116]), .CLK(clk), .RST(rst), .I(g_init[116]), 
        .Q(key[116]) );
  DFF \key_reg[117]  ( .D(nextKey[117]), .CLK(clk), .RST(rst), .I(g_init[117]), 
        .Q(key[117]) );
  DFF \key_reg[118]  ( .D(nextKey[118]), .CLK(clk), .RST(rst), .I(g_init[118]), 
        .Q(key[118]) );
  DFF \key_reg[119]  ( .D(nextKey[119]), .CLK(clk), .RST(rst), .I(g_init[119]), 
        .Q(key[119]) );
  DFF \key_reg[120]  ( .D(nextKey[120]), .CLK(clk), .RST(rst), .I(g_init[120]), 
        .Q(key[120]) );
  DFF \key_reg[121]  ( .D(nextKey[121]), .CLK(clk), .RST(rst), .I(g_init[121]), 
        .Q(key[121]) );
  DFF \key_reg[122]  ( .D(nextKey[122]), .CLK(clk), .RST(rst), .I(g_init[122]), 
        .Q(key[122]) );
  DFF \key_reg[123]  ( .D(nextKey[123]), .CLK(clk), .RST(rst), .I(g_init[123]), 
        .Q(key[123]) );
  DFF \key_reg[124]  ( .D(nextKey[124]), .CLK(clk), .RST(rst), .I(g_init[124]), 
        .Q(key[124]) );
  DFF \key_reg[125]  ( .D(nextKey[125]), .CLK(clk), .RST(rst), .I(g_init[125]), 
        .Q(key[125]) );
  DFF \key_reg[126]  ( .D(nextKey[126]), .CLK(clk), .RST(rst), .I(g_init[126]), 
        .Q(key[126]) );
  DFF \key_reg[127]  ( .D(nextKey[127]), .CLK(clk), .RST(rst), .I(g_init[127]), 
        .Q(key[127]) );
  DFF \msg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(e_init[0]), .Q(msg[0])
         );
  DFF \msg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(e_init[1]), .Q(msg[1])
         );
  DFF \msg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(e_init[2]), .Q(msg[2])
         );
  DFF \msg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(e_init[3]), .Q(msg[3])
         );
  DFF \msg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(e_init[4]), .Q(msg[4])
         );
  DFF \msg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(e_init[5]), .Q(msg[5])
         );
  DFF \msg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(e_init[6]), .Q(msg[6])
         );
  DFF \msg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(e_init[7]), .Q(msg[7])
         );
  DFF \msg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(e_init[8]), .Q(msg[8])
         );
  DFF \msg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(e_init[9]), .Q(msg[9])
         );
  DFF \msg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(e_init[10]), .Q(
        msg[10]) );
  DFF \msg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(e_init[11]), .Q(
        msg[11]) );
  DFF \msg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(e_init[12]), .Q(
        msg[12]) );
  DFF \msg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(e_init[13]), .Q(
        msg[13]) );
  DFF \msg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(e_init[14]), .Q(
        msg[14]) );
  DFF \msg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(e_init[15]), .Q(
        msg[15]) );
  DFF \msg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .I(e_init[16]), .Q(
        msg[16]) );
  DFF \msg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .I(e_init[17]), .Q(
        msg[17]) );
  DFF \msg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .I(e_init[18]), .Q(
        msg[18]) );
  DFF \msg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .I(e_init[19]), .Q(
        msg[19]) );
  DFF \msg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .I(e_init[20]), .Q(
        msg[20]) );
  DFF \msg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .I(e_init[21]), .Q(
        msg[21]) );
  DFF \msg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .I(e_init[22]), .Q(
        msg[22]) );
  DFF \msg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .I(e_init[23]), .Q(
        msg[23]) );
  DFF \msg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .I(e_init[24]), .Q(
        msg[24]) );
  DFF \msg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .I(e_init[25]), .Q(
        msg[25]) );
  DFF \msg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .I(e_init[26]), .Q(
        msg[26]) );
  DFF \msg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .I(e_init[27]), .Q(
        msg[27]) );
  DFF \msg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .I(e_init[28]), .Q(
        msg[28]) );
  DFF \msg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .I(e_init[29]), .Q(
        msg[29]) );
  DFF \msg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .I(e_init[30]), .Q(
        msg[30]) );
  DFF \msg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .I(e_init[31]), .Q(
        msg[31]) );
  DFF \msg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(rst), .I(e_init[32]), .Q(
        msg[32]) );
  DFF \msg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(rst), .I(e_init[33]), .Q(
        msg[33]) );
  DFF \msg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(rst), .I(e_init[34]), .Q(
        msg[34]) );
  DFF \msg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(rst), .I(e_init[35]), .Q(
        msg[35]) );
  DFF \msg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(rst), .I(e_init[36]), .Q(
        msg[36]) );
  DFF \msg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(rst), .I(e_init[37]), .Q(
        msg[37]) );
  DFF \msg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(rst), .I(e_init[38]), .Q(
        msg[38]) );
  DFF \msg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(rst), .I(e_init[39]), .Q(
        msg[39]) );
  DFF \msg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(rst), .I(e_init[40]), .Q(
        msg[40]) );
  DFF \msg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(rst), .I(e_init[41]), .Q(
        msg[41]) );
  DFF \msg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(rst), .I(e_init[42]), .Q(
        msg[42]) );
  DFF \msg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(rst), .I(e_init[43]), .Q(
        msg[43]) );
  DFF \msg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(rst), .I(e_init[44]), .Q(
        msg[44]) );
  DFF \msg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(rst), .I(e_init[45]), .Q(
        msg[45]) );
  DFF \msg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(rst), .I(e_init[46]), .Q(
        msg[46]) );
  DFF \msg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(rst), .I(e_init[47]), .Q(
        msg[47]) );
  DFF \msg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(rst), .I(e_init[48]), .Q(
        msg[48]) );
  DFF \msg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(rst), .I(e_init[49]), .Q(
        msg[49]) );
  DFF \msg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(rst), .I(e_init[50]), .Q(
        msg[50]) );
  DFF \msg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(rst), .I(e_init[51]), .Q(
        msg[51]) );
  DFF \msg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(rst), .I(e_init[52]), .Q(
        msg[52]) );
  DFF \msg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(rst), .I(e_init[53]), .Q(
        msg[53]) );
  DFF \msg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(rst), .I(e_init[54]), .Q(
        msg[54]) );
  DFF \msg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(rst), .I(e_init[55]), .Q(
        msg[55]) );
  DFF \msg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(rst), .I(e_init[56]), .Q(
        msg[56]) );
  DFF \msg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(rst), .I(e_init[57]), .Q(
        msg[57]) );
  DFF \msg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(rst), .I(e_init[58]), .Q(
        msg[58]) );
  DFF \msg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(rst), .I(e_init[59]), .Q(
        msg[59]) );
  DFF \msg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(rst), .I(e_init[60]), .Q(
        msg[60]) );
  DFF \msg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(rst), .I(e_init[61]), .Q(
        msg[61]) );
  DFF \msg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(rst), .I(e_init[62]), .Q(
        msg[62]) );
  DFF \msg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(rst), .I(e_init[63]), .Q(
        msg[63]) );
  DFF \msg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(rst), .I(e_init[64]), .Q(
        msg[64]) );
  DFF \msg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(rst), .I(e_init[65]), .Q(
        msg[65]) );
  DFF \msg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(rst), .I(e_init[66]), .Q(
        msg[66]) );
  DFF \msg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(rst), .I(e_init[67]), .Q(
        msg[67]) );
  DFF \msg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(rst), .I(e_init[68]), .Q(
        msg[68]) );
  DFF \msg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(rst), .I(e_init[69]), .Q(
        msg[69]) );
  DFF \msg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(rst), .I(e_init[70]), .Q(
        msg[70]) );
  DFF \msg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(rst), .I(e_init[71]), .Q(
        msg[71]) );
  DFF \msg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(rst), .I(e_init[72]), .Q(
        msg[72]) );
  DFF \msg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(rst), .I(e_init[73]), .Q(
        msg[73]) );
  DFF \msg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(rst), .I(e_init[74]), .Q(
        msg[74]) );
  DFF \msg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(rst), .I(e_init[75]), .Q(
        msg[75]) );
  DFF \msg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(rst), .I(e_init[76]), .Q(
        msg[76]) );
  DFF \msg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(rst), .I(e_init[77]), .Q(
        msg[77]) );
  DFF \msg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(rst), .I(e_init[78]), .Q(
        msg[78]) );
  DFF \msg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(rst), .I(e_init[79]), .Q(
        msg[79]) );
  DFF \msg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(rst), .I(e_init[80]), .Q(
        msg[80]) );
  DFF \msg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(rst), .I(e_init[81]), .Q(
        msg[81]) );
  DFF \msg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(rst), .I(e_init[82]), .Q(
        msg[82]) );
  DFF \msg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(rst), .I(e_init[83]), .Q(
        msg[83]) );
  DFF \msg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(rst), .I(e_init[84]), .Q(
        msg[84]) );
  DFF \msg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(rst), .I(e_init[85]), .Q(
        msg[85]) );
  DFF \msg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(rst), .I(e_init[86]), .Q(
        msg[86]) );
  DFF \msg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(rst), .I(e_init[87]), .Q(
        msg[87]) );
  DFF \msg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(rst), .I(e_init[88]), .Q(
        msg[88]) );
  DFF \msg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(rst), .I(e_init[89]), .Q(
        msg[89]) );
  DFF \msg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(rst), .I(e_init[90]), .Q(
        msg[90]) );
  DFF \msg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(rst), .I(e_init[91]), .Q(
        msg[91]) );
  DFF \msg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(rst), .I(e_init[92]), .Q(
        msg[92]) );
  DFF \msg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(rst), .I(e_init[93]), .Q(
        msg[93]) );
  DFF \msg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(rst), .I(e_init[94]), .Q(
        msg[94]) );
  DFF \msg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(rst), .I(e_init[95]), .Q(
        msg[95]) );
  DFF \msg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(rst), .I(e_init[96]), .Q(
        msg[96]) );
  DFF \msg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(rst), .I(e_init[97]), .Q(
        msg[97]) );
  DFF \msg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(rst), .I(e_init[98]), .Q(
        msg[98]) );
  DFF \msg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(rst), .I(e_init[99]), .Q(
        msg[99]) );
  DFF \msg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(rst), .I(e_init[100]), .Q(
        msg[100]) );
  DFF \msg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(rst), .I(e_init[101]), .Q(
        msg[101]) );
  DFF \msg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(rst), .I(e_init[102]), .Q(
        msg[102]) );
  DFF \msg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(rst), .I(e_init[103]), .Q(
        msg[103]) );
  DFF \msg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(rst), .I(e_init[104]), .Q(
        msg[104]) );
  DFF \msg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(rst), .I(e_init[105]), .Q(
        msg[105]) );
  DFF \msg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(rst), .I(e_init[106]), .Q(
        msg[106]) );
  DFF \msg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(rst), .I(e_init[107]), .Q(
        msg[107]) );
  DFF \msg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(rst), .I(e_init[108]), .Q(
        msg[108]) );
  DFF \msg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(rst), .I(e_init[109]), .Q(
        msg[109]) );
  DFF \msg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(rst), .I(e_init[110]), .Q(
        msg[110]) );
  DFF \msg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(rst), .I(e_init[111]), .Q(
        msg[111]) );
  DFF \msg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(rst), .I(e_init[112]), .Q(
        msg[112]) );
  DFF \msg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(rst), .I(e_init[113]), .Q(
        msg[113]) );
  DFF \msg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(rst), .I(e_init[114]), .Q(
        msg[114]) );
  DFF \msg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(rst), .I(e_init[115]), .Q(
        msg[115]) );
  DFF \msg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(rst), .I(e_init[116]), .Q(
        msg[116]) );
  DFF \msg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(rst), .I(e_init[117]), .Q(
        msg[117]) );
  DFF \msg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(rst), .I(e_init[118]), .Q(
        msg[118]) );
  DFF \msg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(rst), .I(e_init[119]), .Q(
        msg[119]) );
  DFF \msg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(rst), .I(e_init[120]), .Q(
        msg[120]) );
  DFF \msg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(rst), .I(e_init[121]), .Q(
        msg[121]) );
  DFF \msg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(rst), .I(e_init[122]), .Q(
        msg[122]) );
  DFF \msg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(rst), .I(e_init[123]), .Q(
        msg[123]) );
  DFF \msg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(rst), .I(e_init[124]), .Q(
        msg[124]) );
  DFF \msg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(rst), .I(e_init[125]), .Q(
        msg[125]) );
  DFF \msg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(rst), .I(e_init[126]), .Q(
        msg[126]) );
  DFF \msg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(rst), .I(e_init[127]), .Q(
        msg[127]) );
  XOR \e/U418  ( .A(\e/n180 ), .B(\e/n147 ), .Z(nextKey[0]) );
  XOR \e/U417  ( .A(n544), .B(\e/n188 ), .Z(\e/n147 ) );
  XOR \e/U416  ( .A(\e/n196 ), .B(nextKey[0]), .Z(\e/n260 ) );
  XOR \e/U415  ( .A(\e/n181 ), .B(\e/n148 ), .Z(nextKey[1]) );
  XOR \e/U414  ( .A(n543), .B(\e/n189 ), .Z(\e/n148 ) );
  XOR \e/U413  ( .A(\e/n197 ), .B(nextKey[1]), .Z(\e/n261 ) );
  XOR \e/U412  ( .A(\e/n182 ), .B(\e/n149 ), .Z(nextKey[2]) );
  XOR \e/U411  ( .A(\e/Q[2] ), .B(\e/n190 ), .Z(\e/n149 ) );
  XOR \e/U410  ( .A(\e/n198 ), .B(nextKey[2]), .Z(\e/n262 ) );
  XOR \e/U409  ( .A(\e/n183 ), .B(\e/n150 ), .Z(nextKey[3]) );
  XOR \e/U408  ( .A(\e/Q[3] ), .B(\e/n191 ), .Z(\e/n150 ) );
  XOR \e/U407  ( .A(\e/n199 ), .B(nextKey[3]), .Z(\e/n263 ) );
  XOR \e/U406  ( .A(\e/n184 ), .B(\e/n151 ), .Z(nextKey[4]) );
  XOR \e/U405  ( .A(\e/Q[4] ), .B(\e/n192 ), .Z(\e/n151 ) );
  XOR \e/U404  ( .A(\e/n200 ), .B(nextKey[4]), .Z(\e/n264 ) );
  XOR \e/U403  ( .A(\e/n185 ), .B(\e/n152 ), .Z(nextKey[5]) );
  XOR \e/U402  ( .A(n542), .B(\e/n193 ), .Z(\e/n152 ) );
  XOR \e/U401  ( .A(\e/n201 ), .B(nextKey[5]), .Z(\e/n265 ) );
  XOR \e/U400  ( .A(\e/n186 ), .B(\e/n153 ), .Z(nextKey[6]) );
  XOR \e/U399  ( .A(n541), .B(\e/n194 ), .Z(\e/n153 ) );
  XOR \e/U398  ( .A(\e/n202 ), .B(nextKey[6]), .Z(\e/n266 ) );
  XOR \e/U397  ( .A(\e/n187 ), .B(\e/n154 ), .Z(nextKey[7]) );
  XOR \e/U396  ( .A(\e/Q[7] ), .B(\e/n195 ), .Z(\e/n154 ) );
  XOR \e/U395  ( .A(\e/n203 ), .B(nextKey[7]), .Z(\e/n267 ) );
  XOR \e/U394  ( .A(\e/n98 ), .B(\e/n155 ), .Z(nextKey[40]) );
  XOR \e/U393  ( .A(n540), .B(\e/n204 ), .Z(\e/n155 ) );
  XOR \e/U392  ( .A(\e/n236 ), .B(nextKey[40]), .Z(\e/n268 ) );
  XOR \e/U391  ( .A(\e/n97 ), .B(\e/n156 ), .Z(nextKey[41]) );
  XOR \e/U390  ( .A(n539), .B(\e/n205 ), .Z(\e/n156 ) );
  XOR \e/U389  ( .A(\e/n237 ), .B(nextKey[41]), .Z(\e/n269 ) );
  XOR \e/U388  ( .A(\e/n96 ), .B(\e/n157 ), .Z(nextKey[42]) );
  XOR \e/U387  ( .A(\e/t[10] ), .B(\e/n206 ), .Z(\e/n157 ) );
  XOR \e/U386  ( .A(\e/n238 ), .B(nextKey[42]), .Z(\e/n270 ) );
  XOR \e/U385  ( .A(\e/n95 ), .B(\e/n158 ), .Z(nextKey[43]) );
  XOR \e/U384  ( .A(\e/t[11] ), .B(\e/n207 ), .Z(\e/n158 ) );
  XOR \e/U383  ( .A(\e/n239 ), .B(nextKey[43]), .Z(\e/n271 ) );
  XOR \e/U382  ( .A(\e/n94 ), .B(\e/n159 ), .Z(nextKey[44]) );
  XOR \e/U381  ( .A(\e/t[12] ), .B(\e/n208 ), .Z(\e/n159 ) );
  XOR \e/U380  ( .A(\e/n240 ), .B(nextKey[44]), .Z(\e/n272 ) );
  XOR \e/U379  ( .A(\e/n93 ), .B(\e/n160 ), .Z(nextKey[45]) );
  XOR \e/U378  ( .A(n538), .B(\e/n209 ), .Z(\e/n160 ) );
  XOR \e/U377  ( .A(\e/n241 ), .B(nextKey[45]), .Z(\e/n273 ) );
  XOR \e/U376  ( .A(\e/n92 ), .B(\e/n161 ), .Z(nextKey[46]) );
  XOR \e/U375  ( .A(n537), .B(\e/n210 ), .Z(\e/n161 ) );
  XOR \e/U374  ( .A(\e/n242 ), .B(nextKey[46]), .Z(\e/n274 ) );
  XOR \e/U373  ( .A(\e/n91 ), .B(\e/n162 ), .Z(nextKey[47]) );
  XOR \e/U372  ( .A(\e/t[15] ), .B(\e/n211 ), .Z(\e/n162 ) );
  XOR \e/U371  ( .A(\e/n243 ), .B(nextKey[47]), .Z(\e/n275 ) );
  XOR \e/U370  ( .A(\e/n90 ), .B(\e/n163 ), .Z(nextKey[48]) );
  XOR \e/U369  ( .A(n536), .B(\e/n212 ), .Z(\e/n163 ) );
  XOR \e/U368  ( .A(\e/n244 ), .B(nextKey[48]), .Z(\e/n276 ) );
  XOR \e/U367  ( .A(\e/n89 ), .B(\e/n164 ), .Z(nextKey[49]) );
  XOR \e/U366  ( .A(n535), .B(\e/n213 ), .Z(\e/n164 ) );
  XOR \e/U365  ( .A(\e/n245 ), .B(nextKey[49]), .Z(\e/n277 ) );
  XOR \e/U364  ( .A(\e/n88 ), .B(\e/n165 ), .Z(nextKey[50]) );
  XOR \e/U363  ( .A(\e/t[18] ), .B(\e/n214 ), .Z(\e/n165 ) );
  XOR \e/U362  ( .A(\e/n246 ), .B(nextKey[50]), .Z(\e/n278 ) );
  XOR \e/U361  ( .A(\e/n87 ), .B(\e/n166 ), .Z(nextKey[51]) );
  XOR \e/U360  ( .A(\e/t[19] ), .B(\e/n215 ), .Z(\e/n166 ) );
  XOR \e/U359  ( .A(\e/n247 ), .B(nextKey[51]), .Z(\e/n279 ) );
  XOR \e/U358  ( .A(\e/n86 ), .B(\e/n167 ), .Z(nextKey[52]) );
  XOR \e/U357  ( .A(\e/t[20] ), .B(\e/n216 ), .Z(\e/n167 ) );
  XOR \e/U356  ( .A(\e/n248 ), .B(nextKey[52]), .Z(\e/n280 ) );
  XOR \e/U355  ( .A(\e/n85 ), .B(\e/n168 ), .Z(nextKey[53]) );
  XOR \e/U354  ( .A(n534), .B(\e/n217 ), .Z(\e/n168 ) );
  XOR \e/U353  ( .A(\e/n249 ), .B(nextKey[53]), .Z(\e/n281 ) );
  XOR \e/U352  ( .A(\e/n84 ), .B(\e/n169 ), .Z(nextKey[54]) );
  XOR \e/U351  ( .A(n533), .B(\e/n218 ), .Z(\e/n169 ) );
  XOR \e/U350  ( .A(\e/n250 ), .B(nextKey[54]), .Z(\e/n282 ) );
  XOR \e/U349  ( .A(\e/n83 ), .B(\e/n170 ), .Z(nextKey[55]) );
  XOR \e/U348  ( .A(\e/t[23] ), .B(\e/n219 ), .Z(\e/n170 ) );
  XOR \e/U347  ( .A(\e/n251 ), .B(nextKey[55]), .Z(\e/n283 ) );
  XOR \e/U346  ( .A(\e/n82 ), .B(\e/n171 ), .Z(nextKey[56]) );
  XOR \e/U345  ( .A(n532), .B(\e/n220 ), .Z(\e/n171 ) );
  XOR \e/U344  ( .A(\e/n252 ), .B(nextKey[56]), .Z(\e/n284 ) );
  XOR \e/U343  ( .A(\e/n81 ), .B(\e/n172 ), .Z(nextKey[57]) );
  XOR \e/U342  ( .A(n531), .B(\e/n221 ), .Z(\e/n172 ) );
  XOR \e/U341  ( .A(\e/n253 ), .B(nextKey[57]), .Z(\e/n285 ) );
  XOR \e/U340  ( .A(\e/n80 ), .B(\e/n173 ), .Z(nextKey[58]) );
  XOR \e/U339  ( .A(\e/t[26] ), .B(\e/n222 ), .Z(\e/n173 ) );
  XOR \e/U338  ( .A(\e/n254 ), .B(nextKey[58]), .Z(\e/n286 ) );
  XOR \e/U337  ( .A(\e/n79 ), .B(\e/n174 ), .Z(nextKey[59]) );
  XOR \e/U336  ( .A(\e/t[27] ), .B(\e/n223 ), .Z(\e/n174 ) );
  XOR \e/U335  ( .A(\e/n255 ), .B(nextKey[59]), .Z(\e/n287 ) );
  XOR \e/U334  ( .A(\e/n78 ), .B(\e/n175 ), .Z(nextKey[60]) );
  XOR \e/U333  ( .A(\e/t[28] ), .B(\e/n224 ), .Z(\e/n175 ) );
  XOR \e/U332  ( .A(\e/n256 ), .B(nextKey[60]), .Z(\e/n288 ) );
  XOR \e/U331  ( .A(\e/n77 ), .B(\e/n176 ), .Z(nextKey[61]) );
  XOR \e/U330  ( .A(n530), .B(\e/n225 ), .Z(\e/n176 ) );
  XOR \e/U329  ( .A(\e/n257 ), .B(nextKey[61]), .Z(\e/n289 ) );
  XOR \e/U328  ( .A(\e/n76 ), .B(\e/n177 ), .Z(nextKey[62]) );
  XOR \e/U327  ( .A(n529), .B(\e/n226 ), .Z(\e/n177 ) );
  XOR \e/U326  ( .A(\e/n258 ), .B(nextKey[62]), .Z(\e/n290 ) );
  XOR \e/U325  ( .A(\e/n75 ), .B(\e/n178 ), .Z(nextKey[63]) );
  XOR \e/U324  ( .A(\e/t[31] ), .B(\e/n227 ), .Z(\e/n178 ) );
  XOR \e/U323  ( .A(\e/n259 ), .B(nextKey[63]), .Z(\e/n291 ) );
  XOR \e/U322  ( .A(\e/n228 ), .B(\e/n260 ), .Z(nextKey[64]) );
  XOR \e/U320  ( .A(\e/n229 ), .B(\e/n261 ), .Z(nextKey[65]) );
  XOR \e/U318  ( .A(\e/n230 ), .B(\e/n262 ), .Z(nextKey[66]) );
  XOR \e/U316  ( .A(\e/n231 ), .B(\e/n263 ), .Z(nextKey[67]) );
  XOR \e/U314  ( .A(\e/n232 ), .B(\e/n264 ), .Z(nextKey[68]) );
  XOR \e/U312  ( .A(\e/n233 ), .B(\e/n265 ), .Z(nextKey[69]) );
  XOR \e/U310  ( .A(\e/n234 ), .B(\e/n266 ), .Z(nextKey[70]) );
  XOR \e/U308  ( .A(\e/n235 ), .B(\e/n267 ), .Z(nextKey[71]) );
  XOR \e/U306  ( .A(\e/n66 ), .B(\e/n268 ), .Z(nextKey[104]) );
  XOR \e/U298  ( .A(\e/n58 ), .B(\e/n276 ), .Z(nextKey[112]) );
  XOR \e/U290  ( .A(\e/n50 ), .B(\e/n284 ), .Z(nextKey[120]) );
  XOR \b/SBOX[0].sbox/U157  ( .A(\b/SBOX[0].sbox/z[12] ), .B(
        \b/SBOX[0].sbox/n11 ), .Z(\b/SBOX[0].sbox/n75 ) );
  XOR \b/SBOX[0].sbox/U156  ( .A(\b/SBOX[0].sbox/z[0] ), .B(
        \b/SBOX[0].sbox/z[2] ), .Z(\b/SBOX[0].sbox/n11 ) );
  XOR \b/SBOX[0].sbox/U155  ( .A(\b/SBOX[0].sbox/n13 ), .B(
        \b/SBOX[0].sbox/n12 ), .Z(\b/SBOX[0].sbox/n74 ) );
  XOR \b/SBOX[0].sbox/U154  ( .A(\b/SBOX[0].sbox/z[15] ), .B(
        \b/SBOX[0].sbox/z[16] ), .Z(\b/SBOX[0].sbox/n12 ) );
  XOR \b/SBOX[0].sbox/U153  ( .A(\b/SBOX[0].sbox/z[5] ), .B(
        \b/SBOX[0].sbox/z[13] ), .Z(\b/SBOX[0].sbox/n13 ) );
  XOR \b/SBOX[0].sbox/U152  ( .A(\b/SBOX[0].sbox/n74 ), .B(
        \b/SBOX[0].sbox/n14 ), .Z(\b/SBOX[0].sbox/n88 ) );
  XOR \b/SBOX[0].sbox/U151  ( .A(\b/SBOX[0].sbox/z[3] ), .B(
        \b/SBOX[0].sbox/n75 ), .Z(\b/SBOX[0].sbox/n14 ) );
  XOR \b/SBOX[0].sbox/U150  ( .A(\b/SBOX[0].sbox/n16 ), .B(
        \b/SBOX[0].sbox/n15 ), .Z(\b/SBOX[0].sbox/n89 ) );
  XOR \b/SBOX[0].sbox/U149  ( .A(\b/SBOX[0].sbox/n74 ), .B(
        \b/SBOX[0].sbox/n17 ), .Z(\b/SBOX[0].sbox/n15 ) );
  XOR \b/SBOX[0].sbox/U148  ( .A(\b/SBOX[0].sbox/z[8] ), .B(
        \b/SBOX[0].sbox/z[12] ), .Z(\b/SBOX[0].sbox/n16 ) );
  XOR \b/SBOX[0].sbox/U147  ( .A(\b/SBOX[0].sbox/z[4] ), .B(
        \b/SBOX[0].sbox/z[7] ), .Z(\b/SBOX[0].sbox/n17 ) );
  XOR \b/SBOX[0].sbox/U146  ( .A(\b/SBOX[0].sbox/n75 ), .B(
        \b/SBOX[0].sbox/n18 ), .Z(\b/SBOX[0].sbox/n77 ) );
  XOR \b/SBOX[0].sbox/U145  ( .A(\b/SBOX[0].sbox/z[8] ), .B(
        \b/SBOX[0].sbox/z[14] ), .Z(\b/SBOX[0].sbox/n18 ) );
  XOR \b/SBOX[0].sbox/U144  ( .A(\b/SBOX[0].sbox/n20 ), .B(
        \b/SBOX[0].sbox/n19 ), .Z(\b/SBOX[0].sbox/n90 ) );
  XOR \b/SBOX[0].sbox/U143  ( .A(\b/SBOX[0].sbox/z[17] ), .B(
        \b/SBOX[0].sbox/n77 ), .Z(\b/SBOX[0].sbox/n19 ) );
  XOR \b/SBOX[0].sbox/U142  ( .A(\b/SBOX[0].sbox/z[6] ), .B(
        \b/SBOX[0].sbox/z[15] ), .Z(\b/SBOX[0].sbox/n20 ) );
  XOR \b/SBOX[0].sbox/U141  ( .A(\b/SBOX[0].sbox/z[9] ), .B(
        \b/SBOX[0].sbox/n21 ), .Z(\b/SBOX[0].sbox/n78 ) );
  XOR \b/SBOX[0].sbox/U140  ( .A(\b/SBOX[0].sbox/z[0] ), .B(
        \b/SBOX[0].sbox/z[1] ), .Z(\b/SBOX[0].sbox/n21 ) );
  XOR \b/SBOX[0].sbox/U139  ( .A(\b/SBOX[0].sbox/z[16] ), .B(
        \b/SBOX[0].sbox/n22 ), .Z(\b/SBOX[0].sbox/n76 ) );
  XOR \b/SBOX[0].sbox/U138  ( .A(\b/SBOX[0].sbox/z[10] ), .B(
        \b/SBOX[0].sbox/z[15] ), .Z(\b/SBOX[0].sbox/n22 ) );
  XOR \b/SBOX[0].sbox/U137  ( .A(\b/SBOX[0].sbox/n24 ), .B(
        \b/SBOX[0].sbox/n23 ), .Z(\b/SBOX[0].sbox/n91 ) );
  XOR \b/SBOX[0].sbox/U136  ( .A(\b/SBOX[0].sbox/n78 ), .B(
        \b/SBOX[0].sbox/n76 ), .Z(\b/SBOX[0].sbox/n23 ) );
  XOR \b/SBOX[0].sbox/U135  ( .A(\b/SBOX[0].sbox/z[6] ), .B(
        \b/SBOX[0].sbox/z[7] ), .Z(\b/SBOX[0].sbox/n24 ) );
  XOR \b/SBOX[0].sbox/U134  ( .A(\b/SBOX[0].sbox/z[4] ), .B(
        \b/SBOX[0].sbox/n76 ), .Z(\b/SBOX[0].sbox/n79 ) );
  XOR \b/SBOX[0].sbox/U133  ( .A(\b/SBOX[0].sbox/n79 ), .B(
        \b/SBOX[0].sbox/n25 ), .Z(\b/SBOX[0].sbox/n80 ) );
  XOR \b/SBOX[0].sbox/U132  ( .A(\b/SBOX[0].sbox/z[3] ), .B(
        \b/SBOX[0].sbox/z[7] ), .Z(\b/SBOX[0].sbox/n25 ) );
  XOR \b/SBOX[0].sbox/U131  ( .A(\b/SBOX[0].sbox/n77 ), .B(
        \b/SBOX[0].sbox/n26 ), .Z(shift_row_out[2]) );
  XOR \b/SBOX[0].sbox/U130  ( .A(\b/SBOX[0].sbox/z[11] ), .B(
        \b/SBOX[0].sbox/n80 ), .Z(\b/SBOX[0].sbox/n26 ) );
  XOR \b/SBOX[0].sbox/U129  ( .A(\b/SBOX[0].sbox/n28 ), .B(
        \b/SBOX[0].sbox/n27 ), .Z(shift_row_out[3]) );
  XOR \b/SBOX[0].sbox/U128  ( .A(\b/SBOX[0].sbox/n79 ), .B(
        \b/SBOX[0].sbox/n29 ), .Z(\b/SBOX[0].sbox/n27 ) );
  XOR \b/SBOX[0].sbox/U127  ( .A(\b/SBOX[0].sbox/z[5] ), .B(
        \b/SBOX[0].sbox/z[9] ), .Z(\b/SBOX[0].sbox/n28 ) );
  XOR \b/SBOX[0].sbox/U126  ( .A(\b/SBOX[0].sbox/z[1] ), .B(
        \b/SBOX[0].sbox/z[2] ), .Z(\b/SBOX[0].sbox/n29 ) );
  XOR \b/SBOX[0].sbox/U125  ( .A(\b/SBOX[0].sbox/n78 ), .B(
        \b/SBOX[0].sbox/n30 ), .Z(shift_row_out[4]) );
  XOR \b/SBOX[0].sbox/U124  ( .A(\b/SBOX[0].sbox/z[3] ), .B(
        \b/SBOX[0].sbox/n79 ), .Z(\b/SBOX[0].sbox/n30 ) );
  XOR \b/SBOX[0].sbox/U123  ( .A(\b/SBOX[0].sbox/n80 ), .B(
        \b/SBOX[0].sbox/n31 ), .Z(shift_row_out[7]) );
  XOR \b/SBOX[0].sbox/U122  ( .A(\b/SBOX[0].sbox/z[6] ), .B(
        \b/SBOX[0].sbox/z[9] ), .Z(\b/SBOX[0].sbox/n31 ) );
  XOR \b/SBOX[0].sbox/U121  ( .A(\b/SBOX[0].sbox/n33 ), .B(
        \b/SBOX[0].sbox/n32 ), .Z(\b/SBOX[0].sbox/n81 ) );
  XOR \b/SBOX[0].sbox/U120  ( .A(\b/SBOX[0].sbox/n35 ), .B(
        \b/SBOX[0].sbox/n34 ), .Z(\b/SBOX[0].sbox/n32 ) );
  XOR \b/SBOX[0].sbox/U119  ( .A(msg[5]), .B(msg[1]), .Z(\b/SBOX[0].sbox/n33 )
         );
  XOR \b/SBOX[0].sbox/U118  ( .A(\b/SBOX[0].sbox/t[36] ), .B(
        \b/SBOX[0].sbox/t[39] ), .Z(\b/SBOX[0].sbox/n34 ) );
  XOR \b/SBOX[0].sbox/U117  ( .A(\b/SBOX[0].sbox/t[3] ), .B(
        \b/SBOX[0].sbox/t[8] ), .Z(\b/SBOX[0].sbox/n35 ) );
  XOR \b/SBOX[0].sbox/U116  ( .A(\b/SBOX[0].sbox/n37 ), .B(
        \b/SBOX[0].sbox/n36 ), .Z(\b/SBOX[0].sbox/t[41] ) );
  XOR \b/SBOX[0].sbox/U115  ( .A(\b/SBOX[0].sbox/n81 ), .B(
        \b/SBOX[0].sbox/n38 ), .Z(\b/SBOX[0].sbox/n36 ) );
  XOR \b/SBOX[0].sbox/U114  ( .A(\b/SBOX[0].sbox/t[32] ), .B(msg[7]), .Z(
        \b/SBOX[0].sbox/n37 ) );
  XOR \b/SBOX[0].sbox/U113  ( .A(\b/SBOX[0].sbox/t[5] ), .B(
        \b/SBOX[0].sbox/t[10] ), .Z(\b/SBOX[0].sbox/n38 ) );
  XOR \b/SBOX[0].sbox/U112  ( .A(\b/SBOX[0].sbox/t[2] ), .B(msg[6]), .Z(
        \b/SBOX[0].sbox/n82 ) );
  XOR \b/SBOX[0].sbox/U111  ( .A(\b/SBOX[0].sbox/n40 ), .B(
        \b/SBOX[0].sbox/n39 ), .Z(\b/SBOX[0].sbox/t[45] ) );
  XOR \b/SBOX[0].sbox/U110  ( .A(\b/SBOX[0].sbox/n82 ), .B(
        \b/SBOX[0].sbox/n41 ), .Z(\b/SBOX[0].sbox/n39 ) );
  XOR \b/SBOX[0].sbox/U109  ( .A(msg[4]), .B(\b/SBOX[0].sbox/n81 ), .Z(
        \b/SBOX[0].sbox/n40 ) );
  XOR \b/SBOX[0].sbox/U108  ( .A(\b/SBOX[0].sbox/t[7] ), .B(
        \b/SBOX[0].sbox/t[28] ), .Z(\b/SBOX[0].sbox/n41 ) );
  XOR \b/SBOX[0].sbox/U107  ( .A(\b/SBOX[0].sbox/n82 ), .B(
        \b/SBOX[0].sbox/n42 ), .Z(\b/SBOX[0].sbox/n87 ) );
  XOR \b/SBOX[0].sbox/U106  ( .A(\b/SBOX[0].sbox/t[5] ), .B(msg[4]), .Z(
        \b/SBOX[0].sbox/n42 ) );
  XOR \b/SBOX[0].sbox/U105  ( .A(msg[7]), .B(\b/SBOX[0].sbox/n43 ), .Z(
        \b/SBOX[0].sbox/n83 ) );
  XOR \b/SBOX[0].sbox/U104  ( .A(\b/SBOX[0].sbox/t[7] ), .B(
        \b/SBOX[0].sbox/t[10] ), .Z(\b/SBOX[0].sbox/n43 ) );
  XOR \b/SBOX[0].sbox/U103  ( .A(\b/SBOX[0].sbox/n45 ), .B(
        \b/SBOX[0].sbox/n44 ), .Z(\b/SBOX[0].sbox/t[42] ) );
  XOR \b/SBOX[0].sbox/U102  ( .A(\b/SBOX[0].sbox/n87 ), .B(
        \b/SBOX[0].sbox/n83 ), .Z(\b/SBOX[0].sbox/n44 ) );
  XOR \b/SBOX[0].sbox/U101  ( .A(\b/SBOX[0].sbox/t[28] ), .B(
        \b/SBOX[0].sbox/t[32] ), .Z(\b/SBOX[0].sbox/n45 ) );
  XOR \b/SBOX[0].sbox/U100  ( .A(msg[1]), .B(\b/SBOX[0].sbox/n46 ), .Z(
        \b/SBOX[0].sbox/n85 ) );
  XOR \b/SBOX[0].sbox/U99  ( .A(msg[3]), .B(msg[2]), .Z(\b/SBOX[0].sbox/n46 )
         );
  XOR \b/SBOX[0].sbox/U98  ( .A(msg[5]), .B(\b/SBOX[0].sbox/n85 ), .Z(
        \b/SBOX[0].sbox/y[16] ) );
  XOR \b/SBOX[0].sbox/U97  ( .A(\b/SBOX[0].sbox/y[16] ), .B(
        \b/SBOX[0].sbox/n47 ), .Z(\b/SBOX[0].sbox/n86 ) );
  XOR \b/SBOX[0].sbox/U96  ( .A(\b/SBOX[0].sbox/t[12] ), .B(
        \b/SBOX[0].sbox/t[15] ), .Z(\b/SBOX[0].sbox/n47 ) );
  XOR \b/SBOX[0].sbox/U95  ( .A(\b/SBOX[0].sbox/n86 ), .B(\b/SBOX[0].sbox/n48 ), .Z(\b/SBOX[0].sbox/t[29] ) );
  XOR \b/SBOX[0].sbox/U94  ( .A(\b/SBOX[0].sbox/t[28] ), .B(
        \b/SBOX[0].sbox/n87 ), .Z(\b/SBOX[0].sbox/n48 ) );
  XOR \b/SBOX[0].sbox/U93  ( .A(msg[0]), .B(\b/SBOX[0].sbox/n49 ), .Z(
        \b/SBOX[0].sbox/y[1] ) );
  XOR \b/SBOX[0].sbox/U92  ( .A(msg[6]), .B(msg[5]), .Z(\b/SBOX[0].sbox/n49 )
         );
  XOR \b/SBOX[0].sbox/U91  ( .A(msg[7]), .B(\b/SBOX[0].sbox/y[1] ), .Z(
        \b/SBOX[0].sbox/y[2] ) );
  XOR \b/SBOX[0].sbox/U90  ( .A(\b/SBOX[0].sbox/n51 ), .B(\b/SBOX[0].sbox/n50 ), .Z(\b/SBOX[0].sbox/t[25] ) );
  XOR \b/SBOX[0].sbox/U89  ( .A(\b/SBOX[0].sbox/n53 ), .B(\b/SBOX[0].sbox/n52 ), .Z(\b/SBOX[0].sbox/n50 ) );
  XOR \b/SBOX[0].sbox/U88  ( .A(msg[7]), .B(msg[5]), .Z(\b/SBOX[0].sbox/n51 )
         );
  XOR \b/SBOX[0].sbox/U87  ( .A(\b/SBOX[0].sbox/t[13] ), .B(
        \b/SBOX[0].sbox/t[15] ), .Z(\b/SBOX[0].sbox/n52 ) );
  XOR \b/SBOX[0].sbox/U86  ( .A(\b/SBOX[0].sbox/t[3] ), .B(
        \b/SBOX[0].sbox/t[5] ), .Z(\b/SBOX[0].sbox/n53 ) );
  XOR \b/SBOX[0].sbox/U85  ( .A(\b/SBOX[0].sbox/t[39] ), .B(
        \b/SBOX[0].sbox/t[25] ), .Z(\b/SBOX[0].sbox/t[40] ) );
  XOR \b/SBOX[0].sbox/U84  ( .A(msg[1]), .B(\b/SBOX[0].sbox/y[1] ), .Z(
        \b/SBOX[0].sbox/y[5] ) );
  XOR \b/SBOX[0].sbox/U83  ( .A(\b/SBOX[0].sbox/n55 ), .B(\b/SBOX[0].sbox/n54 ), .Z(\b/SBOX[0].sbox/y[15] ) );
  XOR \b/SBOX[0].sbox/U82  ( .A(msg[3]), .B(msg[1]), .Z(\b/SBOX[0].sbox/n54 )
         );
  XOR \b/SBOX[0].sbox/U81  ( .A(msg[7]), .B(msg[4]), .Z(\b/SBOX[0].sbox/n55 )
         );
  XOR \b/SBOX[0].sbox/U80  ( .A(\b/SBOX[0].sbox/n57 ), .B(\b/SBOX[0].sbox/n56 ), .Z(\b/SBOX[0].sbox/t[21] ) );
  XOR \b/SBOX[0].sbox/U79  ( .A(\b/SBOX[0].sbox/n59 ), .B(\b/SBOX[0].sbox/n58 ), .Z(\b/SBOX[0].sbox/n56 ) );
  XOR \b/SBOX[0].sbox/U78  ( .A(\b/SBOX[0].sbox/y[15] ), .B(
        \b/SBOX[0].sbox/n82 ), .Z(\b/SBOX[0].sbox/n57 ) );
  XOR \b/SBOX[0].sbox/U77  ( .A(\b/SBOX[0].sbox/t[13] ), .B(msg[2]), .Z(
        \b/SBOX[0].sbox/n58 ) );
  XOR \b/SBOX[0].sbox/U76  ( .A(\b/SBOX[0].sbox/t[3] ), .B(
        \b/SBOX[0].sbox/t[12] ), .Z(\b/SBOX[0].sbox/n59 ) );
  XOR \b/SBOX[0].sbox/U75  ( .A(\b/SBOX[0].sbox/t[21] ), .B(
        \b/SBOX[0].sbox/n60 ), .Z(\b/SBOX[0].sbox/t[43] ) );
  XOR \b/SBOX[0].sbox/U74  ( .A(\b/SBOX[0].sbox/t[28] ), .B(
        \b/SBOX[0].sbox/t[39] ), .Z(\b/SBOX[0].sbox/n60 ) );
  XOR \b/SBOX[0].sbox/U73  ( .A(\b/SBOX[0].sbox/n86 ), .B(\b/SBOX[0].sbox/n83 ), .Z(\b/SBOX[0].sbox/t[24] ) );
  XOR \b/SBOX[0].sbox/U72  ( .A(\b/SBOX[0].sbox/t[32] ), .B(
        \b/SBOX[0].sbox/t[24] ), .Z(\b/SBOX[0].sbox/t[33] ) );
  XOR \b/SBOX[0].sbox/U71  ( .A(msg[4]), .B(\b/SBOX[0].sbox/y[1] ), .Z(
        \b/SBOX[0].sbox/y[4] ) );
  XOR \b/SBOX[0].sbox/U70  ( .A(\b/SBOX[0].sbox/n62 ), .B(\b/SBOX[0].sbox/n61 ), .Z(\b/SBOX[0].sbox/t[30] ) );
  XOR \b/SBOX[0].sbox/U69  ( .A(msg[1]), .B(\b/SBOX[0].sbox/n63 ), .Z(
        \b/SBOX[0].sbox/n61 ) );
  XOR \b/SBOX[0].sbox/U68  ( .A(\b/SBOX[0].sbox/t[13] ), .B(
        \b/SBOX[0].sbox/t[15] ), .Z(\b/SBOX[0].sbox/n62 ) );
  XOR \b/SBOX[0].sbox/U67  ( .A(\b/SBOX[0].sbox/t[8] ), .B(
        \b/SBOX[0].sbox/t[10] ), .Z(\b/SBOX[0].sbox/n63 ) );
  XOR \b/SBOX[0].sbox/U66  ( .A(\b/SBOX[0].sbox/t[30] ), .B(
        \b/SBOX[0].sbox/n64 ), .Z(\b/SBOX[0].sbox/t[37] ) );
  XOR \b/SBOX[0].sbox/U65  ( .A(\b/SBOX[0].sbox/t[32] ), .B(
        \b/SBOX[0].sbox/t[36] ), .Z(\b/SBOX[0].sbox/n64 ) );
  XOR \b/SBOX[0].sbox/U64  ( .A(msg[7]), .B(msg[2]), .Z(\b/SBOX[0].sbox/n84 )
         );
  XOR \b/SBOX[0].sbox/U63  ( .A(\b/SBOX[0].sbox/y[5] ), .B(
        \b/SBOX[0].sbox/n84 ), .Z(\b/SBOX[0].sbox/y[3] ) );
  XOR \b/SBOX[0].sbox/U62  ( .A(\b/SBOX[0].sbox/n66 ), .B(\b/SBOX[0].sbox/n65 ), .Z(\b/SBOX[0].sbox/t[23] ) );
  XOR \b/SBOX[0].sbox/U61  ( .A(\b/SBOX[0].sbox/n68 ), .B(\b/SBOX[0].sbox/n67 ), .Z(\b/SBOX[0].sbox/n65 ) );
  XOR \b/SBOX[0].sbox/U60  ( .A(\b/SBOX[0].sbox/n84 ), .B(\b/SBOX[0].sbox/n69 ), .Z(\b/SBOX[0].sbox/n66 ) );
  XOR \b/SBOX[0].sbox/U59  ( .A(msg[5]), .B(msg[3]), .Z(\b/SBOX[0].sbox/n67 )
         );
  XOR \b/SBOX[0].sbox/U58  ( .A(\b/SBOX[0].sbox/t[12] ), .B(
        \b/SBOX[0].sbox/t[13] ), .Z(\b/SBOX[0].sbox/n68 ) );
  XOR \b/SBOX[0].sbox/U57  ( .A(\b/SBOX[0].sbox/t[7] ), .B(
        \b/SBOX[0].sbox/t[8] ), .Z(\b/SBOX[0].sbox/n69 ) );
  XOR \b/SBOX[0].sbox/U56  ( .A(\b/SBOX[0].sbox/t[36] ), .B(
        \b/SBOX[0].sbox/t[23] ), .Z(\b/SBOX[0].sbox/t[44] ) );
  XOR \b/SBOX[0].sbox/U55  ( .A(\b/SBOX[0].sbox/n84 ), .B(\b/SBOX[0].sbox/n70 ), .Z(\b/SBOX[0].sbox/y[12] ) );
  XOR \b/SBOX[0].sbox/U54  ( .A(msg[4]), .B(msg[1]), .Z(\b/SBOX[0].sbox/n70 )
         );
  XOR \b/SBOX[0].sbox/U53  ( .A(\b/SBOX[0].sbox/y[15] ), .B(
        \b/SBOX[0].sbox/n71 ), .Z(\b/SBOX[0].sbox/y[10] ) );
  XOR \b/SBOX[0].sbox/U52  ( .A(msg[6]), .B(msg[5]), .Z(\b/SBOX[0].sbox/n71 )
         );
  XOR \b/SBOX[0].sbox/U51  ( .A(\b/SBOX[0].sbox/n84 ), .B(\b/SBOX[0].sbox/n72 ), .Z(\b/SBOX[0].sbox/y[17] ) );
  XOR \b/SBOX[0].sbox/U50  ( .A(msg[5]), .B(msg[4]), .Z(\b/SBOX[0].sbox/n72 )
         );
  XOR \b/SBOX[0].sbox/U49  ( .A(msg[6]), .B(\b/SBOX[0].sbox/n85 ), .Z(
        \b/SBOX[0].sbox/y[11] ) );
  XOR \b/SBOX[0].sbox/U48  ( .A(msg[0]), .B(\b/SBOX[0].sbox/y[11] ), .Z(
        \b/SBOX[0].sbox/y[7] ) );
  XOR \b/SBOX[0].sbox/U47  ( .A(msg[0]), .B(\b/SBOX[0].sbox/y[15] ), .Z(
        \b/SBOX[0].sbox/y[6] ) );
  XOR \b/SBOX[0].sbox/U46  ( .A(\b/SBOX[0].sbox/t[26] ), .B(
        \b/SBOX[0].sbox/t[24] ), .Z(\b/SBOX[0].sbox/t[27] ) );
  XOR \b/SBOX[0].sbox/U45  ( .A(\b/SBOX[0].sbox/t[36] ), .B(
        \b/SBOX[0].sbox/t[27] ), .Z(\b/SBOX[0].sbox/t[38] ) );
  XOR \b/SBOX[0].sbox/U44  ( .A(\b/SBOX[0].sbox/n86 ), .B(\b/SBOX[0].sbox/n73 ), .Z(\b/SBOX[0].sbox/t[31] ) );
  XOR \b/SBOX[0].sbox/U43  ( .A(\b/SBOX[0].sbox/t[26] ), .B(
        \b/SBOX[0].sbox/n87 ), .Z(\b/SBOX[0].sbox/n73 ) );
  XOR \e/a/SBOX[15].sbox/U157  ( .A(\e/a/SBOX[15].sbox/z[12] ), .B(n3252), .Z(
        n3316) );
  XOR \e/a/SBOX[15].sbox/U156  ( .A(\e/a/SBOX[15].sbox/z[0] ), .B(
        \e/a/SBOX[15].sbox/z[2] ), .Z(n3252) );
  XOR \e/a/SBOX[15].sbox/U155  ( .A(n3254), .B(n3253), .Z(n3315) );
  XOR \e/a/SBOX[15].sbox/U154  ( .A(\e/a/SBOX[15].sbox/z[15] ), .B(
        \e/a/SBOX[15].sbox/z[16] ), .Z(n3253) );
  XOR \e/a/SBOX[15].sbox/U153  ( .A(\e/a/SBOX[15].sbox/z[5] ), .B(
        \e/a/SBOX[15].sbox/z[13] ), .Z(n3254) );
  XOR \e/a/SBOX[15].sbox/U151  ( .A(\e/a/SBOX[15].sbox/z[3] ), .B(n3316), .Z(
        n3255) );
  XOR \e/a/SBOX[15].sbox/U149  ( .A(n3315), .B(n3258), .Z(n3256) );
  XOR \e/a/SBOX[15].sbox/U148  ( .A(\e/a/SBOX[15].sbox/z[8] ), .B(
        \e/a/SBOX[15].sbox/z[12] ), .Z(n3257) );
  XOR \e/a/SBOX[15].sbox/U147  ( .A(\e/a/SBOX[15].sbox/z[4] ), .B(
        \e/a/SBOX[15].sbox/z[7] ), .Z(n3258) );
  XOR \e/a/SBOX[15].sbox/U146  ( .A(n3316), .B(n3259), .Z(n3318) );
  XOR \e/a/SBOX[15].sbox/U145  ( .A(\e/a/SBOX[15].sbox/z[8] ), .B(
        \e/a/SBOX[15].sbox/z[14] ), .Z(n3259) );
  XOR \e/a/SBOX[15].sbox/U143  ( .A(\e/a/SBOX[15].sbox/z[17] ), .B(n3318), .Z(
        n3260) );
  XOR \e/a/SBOX[15].sbox/U142  ( .A(\e/a/SBOX[15].sbox/z[6] ), .B(
        \e/a/SBOX[15].sbox/z[15] ), .Z(n3261) );
  XOR \e/a/SBOX[15].sbox/U141  ( .A(\e/a/SBOX[15].sbox/z[9] ), .B(n3262), .Z(
        n3319) );
  XOR \e/a/SBOX[15].sbox/U140  ( .A(\e/a/SBOX[15].sbox/z[0] ), .B(
        \e/a/SBOX[15].sbox/z[1] ), .Z(n3262) );
  XOR \e/a/SBOX[15].sbox/U139  ( .A(\e/a/SBOX[15].sbox/z[16] ), .B(n3263), .Z(
        n3317) );
  XOR \e/a/SBOX[15].sbox/U138  ( .A(\e/a/SBOX[15].sbox/z[10] ), .B(
        \e/a/SBOX[15].sbox/z[15] ), .Z(n3263) );
  XOR \e/a/SBOX[15].sbox/U136  ( .A(n3319), .B(n3317), .Z(n3264) );
  XOR \e/a/SBOX[15].sbox/U135  ( .A(\e/a/SBOX[15].sbox/z[6] ), .B(
        \e/a/SBOX[15].sbox/z[7] ), .Z(n3265) );
  XOR \e/a/SBOX[15].sbox/U134  ( .A(\e/a/SBOX[15].sbox/z[4] ), .B(n3317), .Z(
        n3320) );
  XOR \e/a/SBOX[15].sbox/U133  ( .A(n3320), .B(n3266), .Z(n3321) );
  XOR \e/a/SBOX[15].sbox/U132  ( .A(\e/a/SBOX[15].sbox/z[3] ), .B(
        \e/a/SBOX[15].sbox/z[7] ), .Z(n3266) );
  XOR \e/a/SBOX[15].sbox/U131  ( .A(n3318), .B(n3267), .Z(\e/t[26] ) );
  XOR \e/a/SBOX[15].sbox/U130  ( .A(\e/a/SBOX[15].sbox/z[11] ), .B(n3321), .Z(
        n3267) );
  XOR \e/a/SBOX[15].sbox/U129  ( .A(n3269), .B(n3268), .Z(\e/t[27] ) );
  XOR \e/a/SBOX[15].sbox/U128  ( .A(n3320), .B(n3270), .Z(n3268) );
  XOR \e/a/SBOX[15].sbox/U127  ( .A(\e/a/SBOX[15].sbox/z[5] ), .B(
        \e/a/SBOX[15].sbox/z[9] ), .Z(n3269) );
  XOR \e/a/SBOX[15].sbox/U126  ( .A(\e/a/SBOX[15].sbox/z[1] ), .B(
        \e/a/SBOX[15].sbox/z[2] ), .Z(n3270) );
  XOR \e/a/SBOX[15].sbox/U125  ( .A(n3319), .B(n3271), .Z(\e/t[28] ) );
  XOR \e/a/SBOX[15].sbox/U124  ( .A(\e/a/SBOX[15].sbox/z[3] ), .B(n3320), .Z(
        n3271) );
  XOR \e/a/SBOX[15].sbox/U123  ( .A(n3321), .B(n3272), .Z(\e/t[31] ) );
  XOR \e/a/SBOX[15].sbox/U122  ( .A(\e/a/SBOX[15].sbox/z[6] ), .B(
        \e/a/SBOX[15].sbox/z[9] ), .Z(n3272) );
  XOR \e/a/SBOX[15].sbox/U121  ( .A(n3274), .B(n3273), .Z(n3322) );
  XOR \e/a/SBOX[15].sbox/U120  ( .A(n3276), .B(n3275), .Z(n3273) );
  XOR \e/a/SBOX[15].sbox/U119  ( .A(\e/w[3][5] ), .B(\e/w[3][1] ), .Z(n3274)
         );
  XOR \e/a/SBOX[15].sbox/U118  ( .A(\e/a/SBOX[15].sbox/t[36] ), .B(
        \e/a/SBOX[15].sbox/t[39] ), .Z(n3275) );
  XOR \e/a/SBOX[15].sbox/U117  ( .A(\e/a/SBOX[15].sbox/t[3] ), .B(
        \e/a/SBOX[15].sbox/t[8] ), .Z(n3276) );
  XOR \e/a/SBOX[15].sbox/U116  ( .A(n3278), .B(n3277), .Z(
        \e/a/SBOX[15].sbox/t[41] ) );
  XOR \e/a/SBOX[15].sbox/U115  ( .A(n3322), .B(n3279), .Z(n3277) );
  XOR \e/a/SBOX[15].sbox/U114  ( .A(\e/a/SBOX[15].sbox/t[32] ), .B(\e/w[3][7] ), .Z(n3278) );
  XOR \e/a/SBOX[15].sbox/U113  ( .A(\e/a/SBOX[15].sbox/t[5] ), .B(
        \e/a/SBOX[15].sbox/t[10] ), .Z(n3279) );
  XOR \e/a/SBOX[15].sbox/U112  ( .A(\e/a/SBOX[15].sbox/t[2] ), .B(\e/w[3][6] ), 
        .Z(n3323) );
  XOR \e/a/SBOX[15].sbox/U111  ( .A(n3281), .B(n3280), .Z(
        \e/a/SBOX[15].sbox/t[45] ) );
  XOR \e/a/SBOX[15].sbox/U110  ( .A(n3323), .B(n3282), .Z(n3280) );
  XOR \e/a/SBOX[15].sbox/U109  ( .A(\e/w[3][4] ), .B(n3322), .Z(n3281) );
  XOR \e/a/SBOX[15].sbox/U108  ( .A(\e/a/SBOX[15].sbox/t[7] ), .B(
        \e/a/SBOX[15].sbox/t[28] ), .Z(n3282) );
  XOR \e/a/SBOX[15].sbox/U107  ( .A(n3323), .B(n3283), .Z(n3328) );
  XOR \e/a/SBOX[15].sbox/U106  ( .A(\e/a/SBOX[15].sbox/t[5] ), .B(\e/w[3][4] ), 
        .Z(n3283) );
  XOR \e/a/SBOX[15].sbox/U105  ( .A(\e/w[3][7] ), .B(n3284), .Z(n3324) );
  XOR \e/a/SBOX[15].sbox/U104  ( .A(\e/a/SBOX[15].sbox/t[7] ), .B(
        \e/a/SBOX[15].sbox/t[10] ), .Z(n3284) );
  XOR \e/a/SBOX[15].sbox/U103  ( .A(n3286), .B(n3285), .Z(
        \e/a/SBOX[15].sbox/t[42] ) );
  XOR \e/a/SBOX[15].sbox/U102  ( .A(n3328), .B(n3324), .Z(n3285) );
  XOR \e/a/SBOX[15].sbox/U101  ( .A(\e/a/SBOX[15].sbox/t[28] ), .B(
        \e/a/SBOX[15].sbox/t[32] ), .Z(n3286) );
  XOR \e/a/SBOX[15].sbox/U100  ( .A(\e/w[3][1] ), .B(n3287), .Z(n3326) );
  XOR \e/a/SBOX[15].sbox/U99  ( .A(\e/w[3][3] ), .B(\e/w[3][2] ), .Z(n3287) );
  XOR \e/a/SBOX[15].sbox/U98  ( .A(\e/w[3][5] ), .B(n3326), .Z(
        \e/a/SBOX[15].sbox/y[16] ) );
  XOR \e/a/SBOX[15].sbox/U97  ( .A(\e/a/SBOX[15].sbox/y[16] ), .B(n3288), .Z(
        n3327) );
  XOR \e/a/SBOX[15].sbox/U96  ( .A(\e/a/SBOX[15].sbox/t[12] ), .B(
        \e/a/SBOX[15].sbox/t[15] ), .Z(n3288) );
  XOR \e/a/SBOX[15].sbox/U95  ( .A(n3327), .B(n3289), .Z(
        \e/a/SBOX[15].sbox/t[29] ) );
  XOR \e/a/SBOX[15].sbox/U94  ( .A(\e/a/SBOX[15].sbox/t[28] ), .B(n3328), .Z(
        n3289) );
  XOR \e/a/SBOX[15].sbox/U93  ( .A(\e/w[3][0] ), .B(n3290), .Z(
        \e/a/SBOX[15].sbox/y[1] ) );
  XOR \e/a/SBOX[15].sbox/U92  ( .A(\e/w[3][6] ), .B(\e/w[3][5] ), .Z(n3290) );
  XOR \e/a/SBOX[15].sbox/U91  ( .A(\e/w[3][7] ), .B(\e/a/SBOX[15].sbox/y[1] ), 
        .Z(\e/a/SBOX[15].sbox/y[2] ) );
  XOR \e/a/SBOX[15].sbox/U90  ( .A(n3292), .B(n3291), .Z(
        \e/a/SBOX[15].sbox/t[25] ) );
  XOR \e/a/SBOX[15].sbox/U89  ( .A(n3294), .B(n3293), .Z(n3291) );
  XOR \e/a/SBOX[15].sbox/U88  ( .A(\e/w[3][7] ), .B(\e/w[3][5] ), .Z(n3292) );
  XOR \e/a/SBOX[15].sbox/U87  ( .A(\e/a/SBOX[15].sbox/t[13] ), .B(
        \e/a/SBOX[15].sbox/t[15] ), .Z(n3293) );
  XOR \e/a/SBOX[15].sbox/U86  ( .A(\e/a/SBOX[15].sbox/t[3] ), .B(
        \e/a/SBOX[15].sbox/t[5] ), .Z(n3294) );
  XOR \e/a/SBOX[15].sbox/U85  ( .A(\e/a/SBOX[15].sbox/t[39] ), .B(
        \e/a/SBOX[15].sbox/t[25] ), .Z(\e/a/SBOX[15].sbox/t[40] ) );
  XOR \e/a/SBOX[15].sbox/U84  ( .A(\e/w[3][1] ), .B(\e/a/SBOX[15].sbox/y[1] ), 
        .Z(\e/a/SBOX[15].sbox/y[5] ) );
  XOR \e/a/SBOX[15].sbox/U83  ( .A(n3296), .B(n3295), .Z(
        \e/a/SBOX[15].sbox/y[15] ) );
  XOR \e/a/SBOX[15].sbox/U82  ( .A(\e/w[3][3] ), .B(\e/w[3][1] ), .Z(n3295) );
  XOR \e/a/SBOX[15].sbox/U81  ( .A(\e/w[3][7] ), .B(\e/w[3][4] ), .Z(n3296) );
  XOR \e/a/SBOX[15].sbox/U80  ( .A(n3298), .B(n3297), .Z(
        \e/a/SBOX[15].sbox/t[21] ) );
  XOR \e/a/SBOX[15].sbox/U79  ( .A(n3300), .B(n3299), .Z(n3297) );
  XOR \e/a/SBOX[15].sbox/U78  ( .A(\e/a/SBOX[15].sbox/y[15] ), .B(n3323), .Z(
        n3298) );
  XOR \e/a/SBOX[15].sbox/U77  ( .A(\e/a/SBOX[15].sbox/t[13] ), .B(\e/w[3][2] ), 
        .Z(n3299) );
  XOR \e/a/SBOX[15].sbox/U76  ( .A(\e/a/SBOX[15].sbox/t[3] ), .B(
        \e/a/SBOX[15].sbox/t[12] ), .Z(n3300) );
  XOR \e/a/SBOX[15].sbox/U75  ( .A(\e/a/SBOX[15].sbox/t[21] ), .B(n3301), .Z(
        \e/a/SBOX[15].sbox/t[43] ) );
  XOR \e/a/SBOX[15].sbox/U74  ( .A(\e/a/SBOX[15].sbox/t[28] ), .B(
        \e/a/SBOX[15].sbox/t[39] ), .Z(n3301) );
  XOR \e/a/SBOX[15].sbox/U73  ( .A(n3327), .B(n3324), .Z(
        \e/a/SBOX[15].sbox/t[24] ) );
  XOR \e/a/SBOX[15].sbox/U72  ( .A(\e/a/SBOX[15].sbox/t[32] ), .B(
        \e/a/SBOX[15].sbox/t[24] ), .Z(\e/a/SBOX[15].sbox/t[33] ) );
  XOR \e/a/SBOX[15].sbox/U71  ( .A(\e/w[3][4] ), .B(\e/a/SBOX[15].sbox/y[1] ), 
        .Z(\e/a/SBOX[15].sbox/y[4] ) );
  XOR \e/a/SBOX[15].sbox/U70  ( .A(n3303), .B(n3302), .Z(
        \e/a/SBOX[15].sbox/t[30] ) );
  XOR \e/a/SBOX[15].sbox/U69  ( .A(\e/w[3][1] ), .B(n3304), .Z(n3302) );
  XOR \e/a/SBOX[15].sbox/U68  ( .A(\e/a/SBOX[15].sbox/t[13] ), .B(
        \e/a/SBOX[15].sbox/t[15] ), .Z(n3303) );
  XOR \e/a/SBOX[15].sbox/U67  ( .A(\e/a/SBOX[15].sbox/t[8] ), .B(
        \e/a/SBOX[15].sbox/t[10] ), .Z(n3304) );
  XOR \e/a/SBOX[15].sbox/U66  ( .A(\e/a/SBOX[15].sbox/t[30] ), .B(n3305), .Z(
        \e/a/SBOX[15].sbox/t[37] ) );
  XOR \e/a/SBOX[15].sbox/U65  ( .A(\e/a/SBOX[15].sbox/t[32] ), .B(
        \e/a/SBOX[15].sbox/t[36] ), .Z(n3305) );
  XOR \e/a/SBOX[15].sbox/U64  ( .A(\e/w[3][7] ), .B(\e/w[3][2] ), .Z(n3325) );
  XOR \e/a/SBOX[15].sbox/U63  ( .A(\e/a/SBOX[15].sbox/y[5] ), .B(n3325), .Z(
        \e/a/SBOX[15].sbox/y[3] ) );
  XOR \e/a/SBOX[15].sbox/U62  ( .A(n3307), .B(n3306), .Z(
        \e/a/SBOX[15].sbox/t[23] ) );
  XOR \e/a/SBOX[15].sbox/U61  ( .A(n3309), .B(n3308), .Z(n3306) );
  XOR \e/a/SBOX[15].sbox/U60  ( .A(n3325), .B(n3310), .Z(n3307) );
  XOR \e/a/SBOX[15].sbox/U59  ( .A(\e/w[3][5] ), .B(\e/w[3][3] ), .Z(n3308) );
  XOR \e/a/SBOX[15].sbox/U58  ( .A(\e/a/SBOX[15].sbox/t[12] ), .B(
        \e/a/SBOX[15].sbox/t[13] ), .Z(n3309) );
  XOR \e/a/SBOX[15].sbox/U57  ( .A(\e/a/SBOX[15].sbox/t[7] ), .B(
        \e/a/SBOX[15].sbox/t[8] ), .Z(n3310) );
  XOR \e/a/SBOX[15].sbox/U56  ( .A(\e/a/SBOX[15].sbox/t[36] ), .B(
        \e/a/SBOX[15].sbox/t[23] ), .Z(\e/a/SBOX[15].sbox/t[44] ) );
  XOR \e/a/SBOX[15].sbox/U55  ( .A(n3325), .B(n3311), .Z(
        \e/a/SBOX[15].sbox/y[12] ) );
  XOR \e/a/SBOX[15].sbox/U54  ( .A(\e/w[3][4] ), .B(\e/w[3][1] ), .Z(n3311) );
  XOR \e/a/SBOX[15].sbox/U53  ( .A(\e/a/SBOX[15].sbox/y[15] ), .B(n3312), .Z(
        \e/a/SBOX[15].sbox/y[10] ) );
  XOR \e/a/SBOX[15].sbox/U52  ( .A(\e/w[3][6] ), .B(\e/w[3][5] ), .Z(n3312) );
  XOR \e/a/SBOX[15].sbox/U51  ( .A(n3325), .B(n3313), .Z(
        \e/a/SBOX[15].sbox/y[17] ) );
  XOR \e/a/SBOX[15].sbox/U50  ( .A(\e/w[3][5] ), .B(\e/w[3][4] ), .Z(n3313) );
  XOR \e/a/SBOX[15].sbox/U49  ( .A(\e/w[3][6] ), .B(n3326), .Z(
        \e/a/SBOX[15].sbox/y[11] ) );
  XOR \e/a/SBOX[15].sbox/U48  ( .A(\e/w[3][0] ), .B(\e/a/SBOX[15].sbox/y[11] ), 
        .Z(\e/a/SBOX[15].sbox/y[7] ) );
  XOR \e/a/SBOX[15].sbox/U47  ( .A(\e/w[3][0] ), .B(\e/a/SBOX[15].sbox/y[15] ), 
        .Z(\e/a/SBOX[15].sbox/y[6] ) );
  XOR \e/a/SBOX[15].sbox/U46  ( .A(\e/a/SBOX[15].sbox/t[26] ), .B(
        \e/a/SBOX[15].sbox/t[24] ), .Z(\e/a/SBOX[15].sbox/t[27] ) );
  XOR \e/a/SBOX[15].sbox/U45  ( .A(\e/a/SBOX[15].sbox/t[36] ), .B(
        \e/a/SBOX[15].sbox/t[27] ), .Z(\e/a/SBOX[15].sbox/t[38] ) );
  XOR \e/a/SBOX[15].sbox/U44  ( .A(n3327), .B(n3314), .Z(
        \e/a/SBOX[15].sbox/t[31] ) );
  XOR \e/a/SBOX[15].sbox/U43  ( .A(\e/a/SBOX[15].sbox/t[26] ), .B(n3328), .Z(
        n3314) );
  XOR \e/a/SBOX[14].sbox/U157  ( .A(\e/a/SBOX[14].sbox/z[12] ), .B(n3175), .Z(
        n3239) );
  XOR \e/a/SBOX[14].sbox/U156  ( .A(\e/a/SBOX[14].sbox/z[0] ), .B(
        \e/a/SBOX[14].sbox/z[2] ), .Z(n3175) );
  XOR \e/a/SBOX[14].sbox/U155  ( .A(n3177), .B(n3176), .Z(n3238) );
  XOR \e/a/SBOX[14].sbox/U154  ( .A(\e/a/SBOX[14].sbox/z[15] ), .B(
        \e/a/SBOX[14].sbox/z[16] ), .Z(n3176) );
  XOR \e/a/SBOX[14].sbox/U153  ( .A(\e/a/SBOX[14].sbox/z[5] ), .B(
        \e/a/SBOX[14].sbox/z[13] ), .Z(n3177) );
  XOR \e/a/SBOX[14].sbox/U151  ( .A(\e/a/SBOX[14].sbox/z[3] ), .B(n3239), .Z(
        n3178) );
  XOR \e/a/SBOX[14].sbox/U149  ( .A(n3238), .B(n3181), .Z(n3179) );
  XOR \e/a/SBOX[14].sbox/U148  ( .A(\e/a/SBOX[14].sbox/z[8] ), .B(
        \e/a/SBOX[14].sbox/z[12] ), .Z(n3180) );
  XOR \e/a/SBOX[14].sbox/U147  ( .A(\e/a/SBOX[14].sbox/z[4] ), .B(
        \e/a/SBOX[14].sbox/z[7] ), .Z(n3181) );
  XOR \e/a/SBOX[14].sbox/U146  ( .A(n3239), .B(n3182), .Z(n3241) );
  XOR \e/a/SBOX[14].sbox/U145  ( .A(\e/a/SBOX[14].sbox/z[8] ), .B(
        \e/a/SBOX[14].sbox/z[14] ), .Z(n3182) );
  XOR \e/a/SBOX[14].sbox/U143  ( .A(\e/a/SBOX[14].sbox/z[17] ), .B(n3241), .Z(
        n3183) );
  XOR \e/a/SBOX[14].sbox/U142  ( .A(\e/a/SBOX[14].sbox/z[6] ), .B(
        \e/a/SBOX[14].sbox/z[15] ), .Z(n3184) );
  XOR \e/a/SBOX[14].sbox/U141  ( .A(\e/a/SBOX[14].sbox/z[9] ), .B(n3185), .Z(
        n3242) );
  XOR \e/a/SBOX[14].sbox/U140  ( .A(\e/a/SBOX[14].sbox/z[0] ), .B(
        \e/a/SBOX[14].sbox/z[1] ), .Z(n3185) );
  XOR \e/a/SBOX[14].sbox/U139  ( .A(\e/a/SBOX[14].sbox/z[16] ), .B(n3186), .Z(
        n3240) );
  XOR \e/a/SBOX[14].sbox/U138  ( .A(\e/a/SBOX[14].sbox/z[10] ), .B(
        \e/a/SBOX[14].sbox/z[15] ), .Z(n3186) );
  XOR \e/a/SBOX[14].sbox/U136  ( .A(n3242), .B(n3240), .Z(n3187) );
  XOR \e/a/SBOX[14].sbox/U135  ( .A(\e/a/SBOX[14].sbox/z[6] ), .B(
        \e/a/SBOX[14].sbox/z[7] ), .Z(n3188) );
  XOR \e/a/SBOX[14].sbox/U134  ( .A(\e/a/SBOX[14].sbox/z[4] ), .B(n3240), .Z(
        n3243) );
  XOR \e/a/SBOX[14].sbox/U133  ( .A(n3243), .B(n3189), .Z(n3244) );
  XOR \e/a/SBOX[14].sbox/U132  ( .A(\e/a/SBOX[14].sbox/z[3] ), .B(
        \e/a/SBOX[14].sbox/z[7] ), .Z(n3189) );
  XOR \e/a/SBOX[14].sbox/U131  ( .A(n3241), .B(n3190), .Z(\e/t[18] ) );
  XOR \e/a/SBOX[14].sbox/U130  ( .A(\e/a/SBOX[14].sbox/z[11] ), .B(n3244), .Z(
        n3190) );
  XOR \e/a/SBOX[14].sbox/U129  ( .A(n3192), .B(n3191), .Z(\e/t[19] ) );
  XOR \e/a/SBOX[14].sbox/U128  ( .A(n3243), .B(n3193), .Z(n3191) );
  XOR \e/a/SBOX[14].sbox/U127  ( .A(\e/a/SBOX[14].sbox/z[5] ), .B(
        \e/a/SBOX[14].sbox/z[9] ), .Z(n3192) );
  XOR \e/a/SBOX[14].sbox/U126  ( .A(\e/a/SBOX[14].sbox/z[1] ), .B(
        \e/a/SBOX[14].sbox/z[2] ), .Z(n3193) );
  XOR \e/a/SBOX[14].sbox/U125  ( .A(n3242), .B(n3194), .Z(\e/t[20] ) );
  XOR \e/a/SBOX[14].sbox/U124  ( .A(\e/a/SBOX[14].sbox/z[3] ), .B(n3243), .Z(
        n3194) );
  XOR \e/a/SBOX[14].sbox/U123  ( .A(n3244), .B(n3195), .Z(\e/t[23] ) );
  XOR \e/a/SBOX[14].sbox/U122  ( .A(\e/a/SBOX[14].sbox/z[6] ), .B(
        \e/a/SBOX[14].sbox/z[9] ), .Z(n3195) );
  XOR \e/a/SBOX[14].sbox/U121  ( .A(n3197), .B(n3196), .Z(n3245) );
  XOR \e/a/SBOX[14].sbox/U120  ( .A(n3199), .B(n3198), .Z(n3196) );
  XOR \e/a/SBOX[14].sbox/U119  ( .A(\e/w[3][29] ), .B(\e/w[3][25] ), .Z(n3197)
         );
  XOR \e/a/SBOX[14].sbox/U118  ( .A(\e/a/SBOX[14].sbox/t[36] ), .B(
        \e/a/SBOX[14].sbox/t[39] ), .Z(n3198) );
  XOR \e/a/SBOX[14].sbox/U117  ( .A(\e/a/SBOX[14].sbox/t[3] ), .B(
        \e/a/SBOX[14].sbox/t[8] ), .Z(n3199) );
  XOR \e/a/SBOX[14].sbox/U116  ( .A(n3201), .B(n3200), .Z(
        \e/a/SBOX[14].sbox/t[41] ) );
  XOR \e/a/SBOX[14].sbox/U115  ( .A(n3245), .B(n3202), .Z(n3200) );
  XOR \e/a/SBOX[14].sbox/U114  ( .A(\e/a/SBOX[14].sbox/t[32] ), .B(
        \e/w[3][31] ), .Z(n3201) );
  XOR \e/a/SBOX[14].sbox/U113  ( .A(\e/a/SBOX[14].sbox/t[5] ), .B(
        \e/a/SBOX[14].sbox/t[10] ), .Z(n3202) );
  XOR \e/a/SBOX[14].sbox/U112  ( .A(\e/a/SBOX[14].sbox/t[2] ), .B(\e/w[3][30] ), .Z(n3246) );
  XOR \e/a/SBOX[14].sbox/U111  ( .A(n3204), .B(n3203), .Z(
        \e/a/SBOX[14].sbox/t[45] ) );
  XOR \e/a/SBOX[14].sbox/U110  ( .A(n3246), .B(n3205), .Z(n3203) );
  XOR \e/a/SBOX[14].sbox/U109  ( .A(\e/w[3][28] ), .B(n3245), .Z(n3204) );
  XOR \e/a/SBOX[14].sbox/U108  ( .A(\e/a/SBOX[14].sbox/t[7] ), .B(
        \e/a/SBOX[14].sbox/t[28] ), .Z(n3205) );
  XOR \e/a/SBOX[14].sbox/U107  ( .A(n3246), .B(n3206), .Z(n3251) );
  XOR \e/a/SBOX[14].sbox/U106  ( .A(\e/a/SBOX[14].sbox/t[5] ), .B(\e/w[3][28] ), .Z(n3206) );
  XOR \e/a/SBOX[14].sbox/U105  ( .A(\e/w[3][31] ), .B(n3207), .Z(n3247) );
  XOR \e/a/SBOX[14].sbox/U104  ( .A(\e/a/SBOX[14].sbox/t[7] ), .B(
        \e/a/SBOX[14].sbox/t[10] ), .Z(n3207) );
  XOR \e/a/SBOX[14].sbox/U103  ( .A(n3209), .B(n3208), .Z(
        \e/a/SBOX[14].sbox/t[42] ) );
  XOR \e/a/SBOX[14].sbox/U102  ( .A(n3251), .B(n3247), .Z(n3208) );
  XOR \e/a/SBOX[14].sbox/U101  ( .A(\e/a/SBOX[14].sbox/t[28] ), .B(
        \e/a/SBOX[14].sbox/t[32] ), .Z(n3209) );
  XOR \e/a/SBOX[14].sbox/U100  ( .A(\e/w[3][25] ), .B(n3210), .Z(n3249) );
  XOR \e/a/SBOX[14].sbox/U99  ( .A(\e/w[3][27] ), .B(\e/w[3][26] ), .Z(n3210)
         );
  XOR \e/a/SBOX[14].sbox/U98  ( .A(\e/w[3][29] ), .B(n3249), .Z(
        \e/a/SBOX[14].sbox/y[16] ) );
  XOR \e/a/SBOX[14].sbox/U97  ( .A(\e/a/SBOX[14].sbox/y[16] ), .B(n3211), .Z(
        n3250) );
  XOR \e/a/SBOX[14].sbox/U96  ( .A(\e/a/SBOX[14].sbox/t[12] ), .B(
        \e/a/SBOX[14].sbox/t[15] ), .Z(n3211) );
  XOR \e/a/SBOX[14].sbox/U95  ( .A(n3250), .B(n3212), .Z(
        \e/a/SBOX[14].sbox/t[29] ) );
  XOR \e/a/SBOX[14].sbox/U94  ( .A(\e/a/SBOX[14].sbox/t[28] ), .B(n3251), .Z(
        n3212) );
  XOR \e/a/SBOX[14].sbox/U93  ( .A(\e/w[3][24] ), .B(n3213), .Z(
        \e/a/SBOX[14].sbox/y[1] ) );
  XOR \e/a/SBOX[14].sbox/U92  ( .A(\e/w[3][30] ), .B(\e/w[3][29] ), .Z(n3213)
         );
  XOR \e/a/SBOX[14].sbox/U91  ( .A(\e/w[3][31] ), .B(\e/a/SBOX[14].sbox/y[1] ), 
        .Z(\e/a/SBOX[14].sbox/y[2] ) );
  XOR \e/a/SBOX[14].sbox/U90  ( .A(n3215), .B(n3214), .Z(
        \e/a/SBOX[14].sbox/t[25] ) );
  XOR \e/a/SBOX[14].sbox/U89  ( .A(n3217), .B(n3216), .Z(n3214) );
  XOR \e/a/SBOX[14].sbox/U88  ( .A(\e/w[3][31] ), .B(\e/w[3][29] ), .Z(n3215)
         );
  XOR \e/a/SBOX[14].sbox/U87  ( .A(\e/a/SBOX[14].sbox/t[13] ), .B(
        \e/a/SBOX[14].sbox/t[15] ), .Z(n3216) );
  XOR \e/a/SBOX[14].sbox/U86  ( .A(\e/a/SBOX[14].sbox/t[3] ), .B(
        \e/a/SBOX[14].sbox/t[5] ), .Z(n3217) );
  XOR \e/a/SBOX[14].sbox/U85  ( .A(\e/a/SBOX[14].sbox/t[39] ), .B(
        \e/a/SBOX[14].sbox/t[25] ), .Z(\e/a/SBOX[14].sbox/t[40] ) );
  XOR \e/a/SBOX[14].sbox/U84  ( .A(\e/w[3][25] ), .B(\e/a/SBOX[14].sbox/y[1] ), 
        .Z(\e/a/SBOX[14].sbox/y[5] ) );
  XOR \e/a/SBOX[14].sbox/U83  ( .A(n3219), .B(n3218), .Z(
        \e/a/SBOX[14].sbox/y[15] ) );
  XOR \e/a/SBOX[14].sbox/U82  ( .A(\e/w[3][27] ), .B(\e/w[3][25] ), .Z(n3218)
         );
  XOR \e/a/SBOX[14].sbox/U81  ( .A(\e/w[3][31] ), .B(\e/w[3][28] ), .Z(n3219)
         );
  XOR \e/a/SBOX[14].sbox/U80  ( .A(n3221), .B(n3220), .Z(
        \e/a/SBOX[14].sbox/t[21] ) );
  XOR \e/a/SBOX[14].sbox/U79  ( .A(n3223), .B(n3222), .Z(n3220) );
  XOR \e/a/SBOX[14].sbox/U78  ( .A(\e/a/SBOX[14].sbox/y[15] ), .B(n3246), .Z(
        n3221) );
  XOR \e/a/SBOX[14].sbox/U77  ( .A(\e/a/SBOX[14].sbox/t[13] ), .B(\e/w[3][26] ), .Z(n3222) );
  XOR \e/a/SBOX[14].sbox/U76  ( .A(\e/a/SBOX[14].sbox/t[3] ), .B(
        \e/a/SBOX[14].sbox/t[12] ), .Z(n3223) );
  XOR \e/a/SBOX[14].sbox/U75  ( .A(\e/a/SBOX[14].sbox/t[21] ), .B(n3224), .Z(
        \e/a/SBOX[14].sbox/t[43] ) );
  XOR \e/a/SBOX[14].sbox/U74  ( .A(\e/a/SBOX[14].sbox/t[28] ), .B(
        \e/a/SBOX[14].sbox/t[39] ), .Z(n3224) );
  XOR \e/a/SBOX[14].sbox/U73  ( .A(n3250), .B(n3247), .Z(
        \e/a/SBOX[14].sbox/t[24] ) );
  XOR \e/a/SBOX[14].sbox/U72  ( .A(\e/a/SBOX[14].sbox/t[32] ), .B(
        \e/a/SBOX[14].sbox/t[24] ), .Z(\e/a/SBOX[14].sbox/t[33] ) );
  XOR \e/a/SBOX[14].sbox/U71  ( .A(\e/w[3][28] ), .B(\e/a/SBOX[14].sbox/y[1] ), 
        .Z(\e/a/SBOX[14].sbox/y[4] ) );
  XOR \e/a/SBOX[14].sbox/U70  ( .A(n3226), .B(n3225), .Z(
        \e/a/SBOX[14].sbox/t[30] ) );
  XOR \e/a/SBOX[14].sbox/U69  ( .A(\e/w[3][25] ), .B(n3227), .Z(n3225) );
  XOR \e/a/SBOX[14].sbox/U68  ( .A(\e/a/SBOX[14].sbox/t[13] ), .B(
        \e/a/SBOX[14].sbox/t[15] ), .Z(n3226) );
  XOR \e/a/SBOX[14].sbox/U67  ( .A(\e/a/SBOX[14].sbox/t[8] ), .B(
        \e/a/SBOX[14].sbox/t[10] ), .Z(n3227) );
  XOR \e/a/SBOX[14].sbox/U66  ( .A(\e/a/SBOX[14].sbox/t[30] ), .B(n3228), .Z(
        \e/a/SBOX[14].sbox/t[37] ) );
  XOR \e/a/SBOX[14].sbox/U65  ( .A(\e/a/SBOX[14].sbox/t[32] ), .B(
        \e/a/SBOX[14].sbox/t[36] ), .Z(n3228) );
  XOR \e/a/SBOX[14].sbox/U64  ( .A(\e/w[3][31] ), .B(\e/w[3][26] ), .Z(n3248)
         );
  XOR \e/a/SBOX[14].sbox/U63  ( .A(\e/a/SBOX[14].sbox/y[5] ), .B(n3248), .Z(
        \e/a/SBOX[14].sbox/y[3] ) );
  XOR \e/a/SBOX[14].sbox/U62  ( .A(n3230), .B(n3229), .Z(
        \e/a/SBOX[14].sbox/t[23] ) );
  XOR \e/a/SBOX[14].sbox/U61  ( .A(n3232), .B(n3231), .Z(n3229) );
  XOR \e/a/SBOX[14].sbox/U60  ( .A(n3248), .B(n3233), .Z(n3230) );
  XOR \e/a/SBOX[14].sbox/U59  ( .A(\e/w[3][29] ), .B(\e/w[3][27] ), .Z(n3231)
         );
  XOR \e/a/SBOX[14].sbox/U58  ( .A(\e/a/SBOX[14].sbox/t[12] ), .B(
        \e/a/SBOX[14].sbox/t[13] ), .Z(n3232) );
  XOR \e/a/SBOX[14].sbox/U57  ( .A(\e/a/SBOX[14].sbox/t[7] ), .B(
        \e/a/SBOX[14].sbox/t[8] ), .Z(n3233) );
  XOR \e/a/SBOX[14].sbox/U56  ( .A(\e/a/SBOX[14].sbox/t[36] ), .B(
        \e/a/SBOX[14].sbox/t[23] ), .Z(\e/a/SBOX[14].sbox/t[44] ) );
  XOR \e/a/SBOX[14].sbox/U55  ( .A(n3248), .B(n3234), .Z(
        \e/a/SBOX[14].sbox/y[12] ) );
  XOR \e/a/SBOX[14].sbox/U54  ( .A(\e/w[3][28] ), .B(\e/w[3][25] ), .Z(n3234)
         );
  XOR \e/a/SBOX[14].sbox/U53  ( .A(\e/a/SBOX[14].sbox/y[15] ), .B(n3235), .Z(
        \e/a/SBOX[14].sbox/y[10] ) );
  XOR \e/a/SBOX[14].sbox/U52  ( .A(\e/w[3][30] ), .B(\e/w[3][29] ), .Z(n3235)
         );
  XOR \e/a/SBOX[14].sbox/U51  ( .A(n3248), .B(n3236), .Z(
        \e/a/SBOX[14].sbox/y[17] ) );
  XOR \e/a/SBOX[14].sbox/U50  ( .A(\e/w[3][29] ), .B(\e/w[3][28] ), .Z(n3236)
         );
  XOR \e/a/SBOX[14].sbox/U49  ( .A(\e/w[3][30] ), .B(n3249), .Z(
        \e/a/SBOX[14].sbox/y[11] ) );
  XOR \e/a/SBOX[14].sbox/U48  ( .A(\e/w[3][24] ), .B(\e/a/SBOX[14].sbox/y[11] ), .Z(\e/a/SBOX[14].sbox/y[7] ) );
  XOR \e/a/SBOX[14].sbox/U47  ( .A(\e/w[3][24] ), .B(\e/a/SBOX[14].sbox/y[15] ), .Z(\e/a/SBOX[14].sbox/y[6] ) );
  XOR \e/a/SBOX[14].sbox/U46  ( .A(\e/a/SBOX[14].sbox/t[26] ), .B(
        \e/a/SBOX[14].sbox/t[24] ), .Z(\e/a/SBOX[14].sbox/t[27] ) );
  XOR \e/a/SBOX[14].sbox/U45  ( .A(\e/a/SBOX[14].sbox/t[36] ), .B(
        \e/a/SBOX[14].sbox/t[27] ), .Z(\e/a/SBOX[14].sbox/t[38] ) );
  XOR \e/a/SBOX[14].sbox/U44  ( .A(n3250), .B(n3237), .Z(
        \e/a/SBOX[14].sbox/t[31] ) );
  XOR \e/a/SBOX[14].sbox/U43  ( .A(\e/a/SBOX[14].sbox/t[26] ), .B(n3251), .Z(
        n3237) );
  XOR \e/a/SBOX[13].sbox/U157  ( .A(\e/a/SBOX[13].sbox/z[12] ), .B(n3098), .Z(
        n3162) );
  XOR \e/a/SBOX[13].sbox/U156  ( .A(\e/a/SBOX[13].sbox/z[0] ), .B(
        \e/a/SBOX[13].sbox/z[2] ), .Z(n3098) );
  XOR \e/a/SBOX[13].sbox/U155  ( .A(n3100), .B(n3099), .Z(n3161) );
  XOR \e/a/SBOX[13].sbox/U154  ( .A(\e/a/SBOX[13].sbox/z[15] ), .B(
        \e/a/SBOX[13].sbox/z[16] ), .Z(n3099) );
  XOR \e/a/SBOX[13].sbox/U153  ( .A(\e/a/SBOX[13].sbox/z[5] ), .B(
        \e/a/SBOX[13].sbox/z[13] ), .Z(n3100) );
  XOR \e/a/SBOX[13].sbox/U151  ( .A(\e/a/SBOX[13].sbox/z[3] ), .B(n3162), .Z(
        n3101) );
  XOR \e/a/SBOX[13].sbox/U149  ( .A(n3161), .B(n3104), .Z(n3102) );
  XOR \e/a/SBOX[13].sbox/U148  ( .A(\e/a/SBOX[13].sbox/z[8] ), .B(
        \e/a/SBOX[13].sbox/z[12] ), .Z(n3103) );
  XOR \e/a/SBOX[13].sbox/U147  ( .A(\e/a/SBOX[13].sbox/z[4] ), .B(
        \e/a/SBOX[13].sbox/z[7] ), .Z(n3104) );
  XOR \e/a/SBOX[13].sbox/U146  ( .A(n3162), .B(n3105), .Z(n3164) );
  XOR \e/a/SBOX[13].sbox/U145  ( .A(\e/a/SBOX[13].sbox/z[8] ), .B(
        \e/a/SBOX[13].sbox/z[14] ), .Z(n3105) );
  XOR \e/a/SBOX[13].sbox/U143  ( .A(\e/a/SBOX[13].sbox/z[17] ), .B(n3164), .Z(
        n3106) );
  XOR \e/a/SBOX[13].sbox/U142  ( .A(\e/a/SBOX[13].sbox/z[6] ), .B(
        \e/a/SBOX[13].sbox/z[15] ), .Z(n3107) );
  XOR \e/a/SBOX[13].sbox/U141  ( .A(\e/a/SBOX[13].sbox/z[9] ), .B(n3108), .Z(
        n3165) );
  XOR \e/a/SBOX[13].sbox/U140  ( .A(\e/a/SBOX[13].sbox/z[0] ), .B(
        \e/a/SBOX[13].sbox/z[1] ), .Z(n3108) );
  XOR \e/a/SBOX[13].sbox/U139  ( .A(\e/a/SBOX[13].sbox/z[16] ), .B(n3109), .Z(
        n3163) );
  XOR \e/a/SBOX[13].sbox/U138  ( .A(\e/a/SBOX[13].sbox/z[10] ), .B(
        \e/a/SBOX[13].sbox/z[15] ), .Z(n3109) );
  XOR \e/a/SBOX[13].sbox/U136  ( .A(n3165), .B(n3163), .Z(n3110) );
  XOR \e/a/SBOX[13].sbox/U135  ( .A(\e/a/SBOX[13].sbox/z[6] ), .B(
        \e/a/SBOX[13].sbox/z[7] ), .Z(n3111) );
  XOR \e/a/SBOX[13].sbox/U134  ( .A(\e/a/SBOX[13].sbox/z[4] ), .B(n3163), .Z(
        n3166) );
  XOR \e/a/SBOX[13].sbox/U133  ( .A(n3166), .B(n3112), .Z(n3167) );
  XOR \e/a/SBOX[13].sbox/U132  ( .A(\e/a/SBOX[13].sbox/z[3] ), .B(
        \e/a/SBOX[13].sbox/z[7] ), .Z(n3112) );
  XOR \e/a/SBOX[13].sbox/U131  ( .A(n3164), .B(n3113), .Z(\e/t[10] ) );
  XOR \e/a/SBOX[13].sbox/U130  ( .A(\e/a/SBOX[13].sbox/z[11] ), .B(n3167), .Z(
        n3113) );
  XOR \e/a/SBOX[13].sbox/U129  ( .A(n3115), .B(n3114), .Z(\e/t[11] ) );
  XOR \e/a/SBOX[13].sbox/U128  ( .A(n3166), .B(n3116), .Z(n3114) );
  XOR \e/a/SBOX[13].sbox/U127  ( .A(\e/a/SBOX[13].sbox/z[5] ), .B(
        \e/a/SBOX[13].sbox/z[9] ), .Z(n3115) );
  XOR \e/a/SBOX[13].sbox/U126  ( .A(\e/a/SBOX[13].sbox/z[1] ), .B(
        \e/a/SBOX[13].sbox/z[2] ), .Z(n3116) );
  XOR \e/a/SBOX[13].sbox/U125  ( .A(n3165), .B(n3117), .Z(\e/t[12] ) );
  XOR \e/a/SBOX[13].sbox/U124  ( .A(\e/a/SBOX[13].sbox/z[3] ), .B(n3166), .Z(
        n3117) );
  XOR \e/a/SBOX[13].sbox/U123  ( .A(n3167), .B(n3118), .Z(\e/t[15] ) );
  XOR \e/a/SBOX[13].sbox/U122  ( .A(\e/a/SBOX[13].sbox/z[6] ), .B(
        \e/a/SBOX[13].sbox/z[9] ), .Z(n3118) );
  XOR \e/a/SBOX[13].sbox/U121  ( .A(n3120), .B(n3119), .Z(n3168) );
  XOR \e/a/SBOX[13].sbox/U120  ( .A(n3122), .B(n3121), .Z(n3119) );
  XOR \e/a/SBOX[13].sbox/U119  ( .A(\e/w[3][21] ), .B(\e/w[3][17] ), .Z(n3120)
         );
  XOR \e/a/SBOX[13].sbox/U118  ( .A(\e/a/SBOX[13].sbox/t[36] ), .B(
        \e/a/SBOX[13].sbox/t[39] ), .Z(n3121) );
  XOR \e/a/SBOX[13].sbox/U117  ( .A(\e/a/SBOX[13].sbox/t[3] ), .B(
        \e/a/SBOX[13].sbox/t[8] ), .Z(n3122) );
  XOR \e/a/SBOX[13].sbox/U116  ( .A(n3124), .B(n3123), .Z(
        \e/a/SBOX[13].sbox/t[41] ) );
  XOR \e/a/SBOX[13].sbox/U115  ( .A(n3168), .B(n3125), .Z(n3123) );
  XOR \e/a/SBOX[13].sbox/U114  ( .A(\e/a/SBOX[13].sbox/t[32] ), .B(
        \e/w[3][23] ), .Z(n3124) );
  XOR \e/a/SBOX[13].sbox/U113  ( .A(\e/a/SBOX[13].sbox/t[5] ), .B(
        \e/a/SBOX[13].sbox/t[10] ), .Z(n3125) );
  XOR \e/a/SBOX[13].sbox/U112  ( .A(\e/a/SBOX[13].sbox/t[2] ), .B(\e/w[3][22] ), .Z(n3169) );
  XOR \e/a/SBOX[13].sbox/U111  ( .A(n3127), .B(n3126), .Z(
        \e/a/SBOX[13].sbox/t[45] ) );
  XOR \e/a/SBOX[13].sbox/U110  ( .A(n3169), .B(n3128), .Z(n3126) );
  XOR \e/a/SBOX[13].sbox/U109  ( .A(\e/w[3][20] ), .B(n3168), .Z(n3127) );
  XOR \e/a/SBOX[13].sbox/U108  ( .A(\e/a/SBOX[13].sbox/t[7] ), .B(
        \e/a/SBOX[13].sbox/t[28] ), .Z(n3128) );
  XOR \e/a/SBOX[13].sbox/U107  ( .A(n3169), .B(n3129), .Z(n3174) );
  XOR \e/a/SBOX[13].sbox/U106  ( .A(\e/a/SBOX[13].sbox/t[5] ), .B(\e/w[3][20] ), .Z(n3129) );
  XOR \e/a/SBOX[13].sbox/U105  ( .A(\e/w[3][23] ), .B(n3130), .Z(n3170) );
  XOR \e/a/SBOX[13].sbox/U104  ( .A(\e/a/SBOX[13].sbox/t[7] ), .B(
        \e/a/SBOX[13].sbox/t[10] ), .Z(n3130) );
  XOR \e/a/SBOX[13].sbox/U103  ( .A(n3132), .B(n3131), .Z(
        \e/a/SBOX[13].sbox/t[42] ) );
  XOR \e/a/SBOX[13].sbox/U102  ( .A(n3174), .B(n3170), .Z(n3131) );
  XOR \e/a/SBOX[13].sbox/U101  ( .A(\e/a/SBOX[13].sbox/t[28] ), .B(
        \e/a/SBOX[13].sbox/t[32] ), .Z(n3132) );
  XOR \e/a/SBOX[13].sbox/U100  ( .A(\e/w[3][17] ), .B(n3133), .Z(n3172) );
  XOR \e/a/SBOX[13].sbox/U99  ( .A(\e/w[3][19] ), .B(\e/w[3][18] ), .Z(n3133)
         );
  XOR \e/a/SBOX[13].sbox/U98  ( .A(\e/w[3][21] ), .B(n3172), .Z(
        \e/a/SBOX[13].sbox/y[16] ) );
  XOR \e/a/SBOX[13].sbox/U97  ( .A(\e/a/SBOX[13].sbox/y[16] ), .B(n3134), .Z(
        n3173) );
  XOR \e/a/SBOX[13].sbox/U96  ( .A(\e/a/SBOX[13].sbox/t[12] ), .B(
        \e/a/SBOX[13].sbox/t[15] ), .Z(n3134) );
  XOR \e/a/SBOX[13].sbox/U95  ( .A(n3173), .B(n3135), .Z(
        \e/a/SBOX[13].sbox/t[29] ) );
  XOR \e/a/SBOX[13].sbox/U94  ( .A(\e/a/SBOX[13].sbox/t[28] ), .B(n3174), .Z(
        n3135) );
  XOR \e/a/SBOX[13].sbox/U93  ( .A(\e/w[3][16] ), .B(n3136), .Z(
        \e/a/SBOX[13].sbox/y[1] ) );
  XOR \e/a/SBOX[13].sbox/U92  ( .A(\e/w[3][22] ), .B(\e/w[3][21] ), .Z(n3136)
         );
  XOR \e/a/SBOX[13].sbox/U91  ( .A(\e/w[3][23] ), .B(\e/a/SBOX[13].sbox/y[1] ), 
        .Z(\e/a/SBOX[13].sbox/y[2] ) );
  XOR \e/a/SBOX[13].sbox/U90  ( .A(n3138), .B(n3137), .Z(
        \e/a/SBOX[13].sbox/t[25] ) );
  XOR \e/a/SBOX[13].sbox/U89  ( .A(n3140), .B(n3139), .Z(n3137) );
  XOR \e/a/SBOX[13].sbox/U88  ( .A(\e/w[3][23] ), .B(\e/w[3][21] ), .Z(n3138)
         );
  XOR \e/a/SBOX[13].sbox/U87  ( .A(\e/a/SBOX[13].sbox/t[13] ), .B(
        \e/a/SBOX[13].sbox/t[15] ), .Z(n3139) );
  XOR \e/a/SBOX[13].sbox/U86  ( .A(\e/a/SBOX[13].sbox/t[3] ), .B(
        \e/a/SBOX[13].sbox/t[5] ), .Z(n3140) );
  XOR \e/a/SBOX[13].sbox/U85  ( .A(\e/a/SBOX[13].sbox/t[39] ), .B(
        \e/a/SBOX[13].sbox/t[25] ), .Z(\e/a/SBOX[13].sbox/t[40] ) );
  XOR \e/a/SBOX[13].sbox/U84  ( .A(\e/w[3][17] ), .B(\e/a/SBOX[13].sbox/y[1] ), 
        .Z(\e/a/SBOX[13].sbox/y[5] ) );
  XOR \e/a/SBOX[13].sbox/U83  ( .A(n3142), .B(n3141), .Z(
        \e/a/SBOX[13].sbox/y[15] ) );
  XOR \e/a/SBOX[13].sbox/U82  ( .A(\e/w[3][19] ), .B(\e/w[3][17] ), .Z(n3141)
         );
  XOR \e/a/SBOX[13].sbox/U81  ( .A(\e/w[3][23] ), .B(\e/w[3][20] ), .Z(n3142)
         );
  XOR \e/a/SBOX[13].sbox/U80  ( .A(n3144), .B(n3143), .Z(
        \e/a/SBOX[13].sbox/t[21] ) );
  XOR \e/a/SBOX[13].sbox/U79  ( .A(n3146), .B(n3145), .Z(n3143) );
  XOR \e/a/SBOX[13].sbox/U78  ( .A(\e/a/SBOX[13].sbox/y[15] ), .B(n3169), .Z(
        n3144) );
  XOR \e/a/SBOX[13].sbox/U77  ( .A(\e/a/SBOX[13].sbox/t[13] ), .B(\e/w[3][18] ), .Z(n3145) );
  XOR \e/a/SBOX[13].sbox/U76  ( .A(\e/a/SBOX[13].sbox/t[3] ), .B(
        \e/a/SBOX[13].sbox/t[12] ), .Z(n3146) );
  XOR \e/a/SBOX[13].sbox/U75  ( .A(\e/a/SBOX[13].sbox/t[21] ), .B(n3147), .Z(
        \e/a/SBOX[13].sbox/t[43] ) );
  XOR \e/a/SBOX[13].sbox/U74  ( .A(\e/a/SBOX[13].sbox/t[28] ), .B(
        \e/a/SBOX[13].sbox/t[39] ), .Z(n3147) );
  XOR \e/a/SBOX[13].sbox/U73  ( .A(n3173), .B(n3170), .Z(
        \e/a/SBOX[13].sbox/t[24] ) );
  XOR \e/a/SBOX[13].sbox/U72  ( .A(\e/a/SBOX[13].sbox/t[32] ), .B(
        \e/a/SBOX[13].sbox/t[24] ), .Z(\e/a/SBOX[13].sbox/t[33] ) );
  XOR \e/a/SBOX[13].sbox/U71  ( .A(\e/w[3][20] ), .B(\e/a/SBOX[13].sbox/y[1] ), 
        .Z(\e/a/SBOX[13].sbox/y[4] ) );
  XOR \e/a/SBOX[13].sbox/U70  ( .A(n3149), .B(n3148), .Z(
        \e/a/SBOX[13].sbox/t[30] ) );
  XOR \e/a/SBOX[13].sbox/U69  ( .A(\e/w[3][17] ), .B(n3150), .Z(n3148) );
  XOR \e/a/SBOX[13].sbox/U68  ( .A(\e/a/SBOX[13].sbox/t[13] ), .B(
        \e/a/SBOX[13].sbox/t[15] ), .Z(n3149) );
  XOR \e/a/SBOX[13].sbox/U67  ( .A(\e/a/SBOX[13].sbox/t[8] ), .B(
        \e/a/SBOX[13].sbox/t[10] ), .Z(n3150) );
  XOR \e/a/SBOX[13].sbox/U66  ( .A(\e/a/SBOX[13].sbox/t[30] ), .B(n3151), .Z(
        \e/a/SBOX[13].sbox/t[37] ) );
  XOR \e/a/SBOX[13].sbox/U65  ( .A(\e/a/SBOX[13].sbox/t[32] ), .B(
        \e/a/SBOX[13].sbox/t[36] ), .Z(n3151) );
  XOR \e/a/SBOX[13].sbox/U64  ( .A(\e/w[3][23] ), .B(\e/w[3][18] ), .Z(n3171)
         );
  XOR \e/a/SBOX[13].sbox/U63  ( .A(\e/a/SBOX[13].sbox/y[5] ), .B(n3171), .Z(
        \e/a/SBOX[13].sbox/y[3] ) );
  XOR \e/a/SBOX[13].sbox/U62  ( .A(n3153), .B(n3152), .Z(
        \e/a/SBOX[13].sbox/t[23] ) );
  XOR \e/a/SBOX[13].sbox/U61  ( .A(n3155), .B(n3154), .Z(n3152) );
  XOR \e/a/SBOX[13].sbox/U60  ( .A(n3171), .B(n3156), .Z(n3153) );
  XOR \e/a/SBOX[13].sbox/U59  ( .A(\e/w[3][21] ), .B(\e/w[3][19] ), .Z(n3154)
         );
  XOR \e/a/SBOX[13].sbox/U58  ( .A(\e/a/SBOX[13].sbox/t[12] ), .B(
        \e/a/SBOX[13].sbox/t[13] ), .Z(n3155) );
  XOR \e/a/SBOX[13].sbox/U57  ( .A(\e/a/SBOX[13].sbox/t[7] ), .B(
        \e/a/SBOX[13].sbox/t[8] ), .Z(n3156) );
  XOR \e/a/SBOX[13].sbox/U56  ( .A(\e/a/SBOX[13].sbox/t[36] ), .B(
        \e/a/SBOX[13].sbox/t[23] ), .Z(\e/a/SBOX[13].sbox/t[44] ) );
  XOR \e/a/SBOX[13].sbox/U55  ( .A(n3171), .B(n3157), .Z(
        \e/a/SBOX[13].sbox/y[12] ) );
  XOR \e/a/SBOX[13].sbox/U54  ( .A(\e/w[3][20] ), .B(\e/w[3][17] ), .Z(n3157)
         );
  XOR \e/a/SBOX[13].sbox/U53  ( .A(\e/a/SBOX[13].sbox/y[15] ), .B(n3158), .Z(
        \e/a/SBOX[13].sbox/y[10] ) );
  XOR \e/a/SBOX[13].sbox/U52  ( .A(\e/w[3][22] ), .B(\e/w[3][21] ), .Z(n3158)
         );
  XOR \e/a/SBOX[13].sbox/U51  ( .A(n3171), .B(n3159), .Z(
        \e/a/SBOX[13].sbox/y[17] ) );
  XOR \e/a/SBOX[13].sbox/U50  ( .A(\e/w[3][21] ), .B(\e/w[3][20] ), .Z(n3159)
         );
  XOR \e/a/SBOX[13].sbox/U49  ( .A(\e/w[3][22] ), .B(n3172), .Z(
        \e/a/SBOX[13].sbox/y[11] ) );
  XOR \e/a/SBOX[13].sbox/U48  ( .A(\e/w[3][16] ), .B(\e/a/SBOX[13].sbox/y[11] ), .Z(\e/a/SBOX[13].sbox/y[7] ) );
  XOR \e/a/SBOX[13].sbox/U47  ( .A(\e/w[3][16] ), .B(\e/a/SBOX[13].sbox/y[15] ), .Z(\e/a/SBOX[13].sbox/y[6] ) );
  XOR \e/a/SBOX[13].sbox/U46  ( .A(\e/a/SBOX[13].sbox/t[26] ), .B(
        \e/a/SBOX[13].sbox/t[24] ), .Z(\e/a/SBOX[13].sbox/t[27] ) );
  XOR \e/a/SBOX[13].sbox/U45  ( .A(\e/a/SBOX[13].sbox/t[36] ), .B(
        \e/a/SBOX[13].sbox/t[27] ), .Z(\e/a/SBOX[13].sbox/t[38] ) );
  XOR \e/a/SBOX[13].sbox/U44  ( .A(n3173), .B(n3160), .Z(
        \e/a/SBOX[13].sbox/t[31] ) );
  XOR \e/a/SBOX[13].sbox/U43  ( .A(\e/a/SBOX[13].sbox/t[26] ), .B(n3174), .Z(
        n3160) );
  XOR \e/a/SBOX[12].sbox/U157  ( .A(\e/a/SBOX[12].sbox/z[12] ), .B(n3021), .Z(
        n3085) );
  XOR \e/a/SBOX[12].sbox/U156  ( .A(\e/a/SBOX[12].sbox/z[0] ), .B(
        \e/a/SBOX[12].sbox/z[2] ), .Z(n3021) );
  XOR \e/a/SBOX[12].sbox/U155  ( .A(n3023), .B(n3022), .Z(n3084) );
  XOR \e/a/SBOX[12].sbox/U154  ( .A(\e/a/SBOX[12].sbox/z[15] ), .B(
        \e/a/SBOX[12].sbox/z[16] ), .Z(n3022) );
  XOR \e/a/SBOX[12].sbox/U153  ( .A(\e/a/SBOX[12].sbox/z[5] ), .B(
        \e/a/SBOX[12].sbox/z[13] ), .Z(n3023) );
  XOR \e/a/SBOX[12].sbox/U151  ( .A(\e/a/SBOX[12].sbox/z[3] ), .B(n3085), .Z(
        n3024) );
  XOR \e/a/SBOX[12].sbox/U149  ( .A(n3084), .B(n3027), .Z(n3025) );
  XOR \e/a/SBOX[12].sbox/U148  ( .A(\e/a/SBOX[12].sbox/z[8] ), .B(
        \e/a/SBOX[12].sbox/z[12] ), .Z(n3026) );
  XOR \e/a/SBOX[12].sbox/U147  ( .A(\e/a/SBOX[12].sbox/z[4] ), .B(
        \e/a/SBOX[12].sbox/z[7] ), .Z(n3027) );
  XOR \e/a/SBOX[12].sbox/U146  ( .A(n3085), .B(n3028), .Z(n3087) );
  XOR \e/a/SBOX[12].sbox/U145  ( .A(\e/a/SBOX[12].sbox/z[8] ), .B(
        \e/a/SBOX[12].sbox/z[14] ), .Z(n3028) );
  XOR \e/a/SBOX[12].sbox/U143  ( .A(\e/a/SBOX[12].sbox/z[17] ), .B(n3087), .Z(
        n3029) );
  XOR \e/a/SBOX[12].sbox/U142  ( .A(\e/a/SBOX[12].sbox/z[6] ), .B(
        \e/a/SBOX[12].sbox/z[15] ), .Z(n3030) );
  XOR \e/a/SBOX[12].sbox/U141  ( .A(\e/a/SBOX[12].sbox/z[9] ), .B(n3031), .Z(
        n3088) );
  XOR \e/a/SBOX[12].sbox/U140  ( .A(\e/a/SBOX[12].sbox/z[0] ), .B(
        \e/a/SBOX[12].sbox/z[1] ), .Z(n3031) );
  XOR \e/a/SBOX[12].sbox/U139  ( .A(\e/a/SBOX[12].sbox/z[16] ), .B(n3032), .Z(
        n3086) );
  XOR \e/a/SBOX[12].sbox/U138  ( .A(\e/a/SBOX[12].sbox/z[10] ), .B(
        \e/a/SBOX[12].sbox/z[15] ), .Z(n3032) );
  XOR \e/a/SBOX[12].sbox/U136  ( .A(n3088), .B(n3086), .Z(n3033) );
  XOR \e/a/SBOX[12].sbox/U135  ( .A(\e/a/SBOX[12].sbox/z[6] ), .B(
        \e/a/SBOX[12].sbox/z[7] ), .Z(n3034) );
  XOR \e/a/SBOX[12].sbox/U134  ( .A(\e/a/SBOX[12].sbox/z[4] ), .B(n3086), .Z(
        n3089) );
  XOR \e/a/SBOX[12].sbox/U133  ( .A(n3089), .B(n3035), .Z(n3090) );
  XOR \e/a/SBOX[12].sbox/U132  ( .A(\e/a/SBOX[12].sbox/z[3] ), .B(
        \e/a/SBOX[12].sbox/z[7] ), .Z(n3035) );
  XOR \e/a/SBOX[12].sbox/U131  ( .A(n3087), .B(n3036), .Z(\e/Q[2] ) );
  XOR \e/a/SBOX[12].sbox/U130  ( .A(\e/a/SBOX[12].sbox/z[11] ), .B(n3090), .Z(
        n3036) );
  XOR \e/a/SBOX[12].sbox/U129  ( .A(n3038), .B(n3037), .Z(\e/Q[3] ) );
  XOR \e/a/SBOX[12].sbox/U128  ( .A(n3089), .B(n3039), .Z(n3037) );
  XOR \e/a/SBOX[12].sbox/U127  ( .A(\e/a/SBOX[12].sbox/z[5] ), .B(
        \e/a/SBOX[12].sbox/z[9] ), .Z(n3038) );
  XOR \e/a/SBOX[12].sbox/U126  ( .A(\e/a/SBOX[12].sbox/z[1] ), .B(
        \e/a/SBOX[12].sbox/z[2] ), .Z(n3039) );
  XOR \e/a/SBOX[12].sbox/U125  ( .A(n3088), .B(n3040), .Z(\e/Q[4] ) );
  XOR \e/a/SBOX[12].sbox/U124  ( .A(\e/a/SBOX[12].sbox/z[3] ), .B(n3089), .Z(
        n3040) );
  XOR \e/a/SBOX[12].sbox/U123  ( .A(n3090), .B(n3041), .Z(\e/Q[7] ) );
  XOR \e/a/SBOX[12].sbox/U122  ( .A(\e/a/SBOX[12].sbox/z[6] ), .B(
        \e/a/SBOX[12].sbox/z[9] ), .Z(n3041) );
  XOR \e/a/SBOX[12].sbox/U121  ( .A(n3043), .B(n3042), .Z(n3091) );
  XOR \e/a/SBOX[12].sbox/U120  ( .A(n3045), .B(n3044), .Z(n3042) );
  XOR \e/a/SBOX[12].sbox/U119  ( .A(\e/w[3][13] ), .B(\e/w[3][9] ), .Z(n3043)
         );
  XOR \e/a/SBOX[12].sbox/U118  ( .A(\e/a/SBOX[12].sbox/t[36] ), .B(
        \e/a/SBOX[12].sbox/t[39] ), .Z(n3044) );
  XOR \e/a/SBOX[12].sbox/U117  ( .A(\e/a/SBOX[12].sbox/t[3] ), .B(
        \e/a/SBOX[12].sbox/t[8] ), .Z(n3045) );
  XOR \e/a/SBOX[12].sbox/U116  ( .A(n3047), .B(n3046), .Z(
        \e/a/SBOX[12].sbox/t[41] ) );
  XOR \e/a/SBOX[12].sbox/U115  ( .A(n3091), .B(n3048), .Z(n3046) );
  XOR \e/a/SBOX[12].sbox/U114  ( .A(\e/a/SBOX[12].sbox/t[32] ), .B(
        \e/w[3][15] ), .Z(n3047) );
  XOR \e/a/SBOX[12].sbox/U113  ( .A(\e/a/SBOX[12].sbox/t[5] ), .B(
        \e/a/SBOX[12].sbox/t[10] ), .Z(n3048) );
  XOR \e/a/SBOX[12].sbox/U112  ( .A(\e/a/SBOX[12].sbox/t[2] ), .B(\e/w[3][14] ), .Z(n3092) );
  XOR \e/a/SBOX[12].sbox/U111  ( .A(n3050), .B(n3049), .Z(
        \e/a/SBOX[12].sbox/t[45] ) );
  XOR \e/a/SBOX[12].sbox/U110  ( .A(n3092), .B(n3051), .Z(n3049) );
  XOR \e/a/SBOX[12].sbox/U109  ( .A(\e/w[3][12] ), .B(n3091), .Z(n3050) );
  XOR \e/a/SBOX[12].sbox/U108  ( .A(\e/a/SBOX[12].sbox/t[7] ), .B(
        \e/a/SBOX[12].sbox/t[28] ), .Z(n3051) );
  XOR \e/a/SBOX[12].sbox/U107  ( .A(n3092), .B(n3052), .Z(n3097) );
  XOR \e/a/SBOX[12].sbox/U106  ( .A(\e/a/SBOX[12].sbox/t[5] ), .B(\e/w[3][12] ), .Z(n3052) );
  XOR \e/a/SBOX[12].sbox/U105  ( .A(\e/w[3][15] ), .B(n3053), .Z(n3093) );
  XOR \e/a/SBOX[12].sbox/U104  ( .A(\e/a/SBOX[12].sbox/t[7] ), .B(
        \e/a/SBOX[12].sbox/t[10] ), .Z(n3053) );
  XOR \e/a/SBOX[12].sbox/U103  ( .A(n3055), .B(n3054), .Z(
        \e/a/SBOX[12].sbox/t[42] ) );
  XOR \e/a/SBOX[12].sbox/U102  ( .A(n3097), .B(n3093), .Z(n3054) );
  XOR \e/a/SBOX[12].sbox/U101  ( .A(\e/a/SBOX[12].sbox/t[28] ), .B(
        \e/a/SBOX[12].sbox/t[32] ), .Z(n3055) );
  XOR \e/a/SBOX[12].sbox/U100  ( .A(\e/w[3][9] ), .B(n3056), .Z(n3095) );
  XOR \e/a/SBOX[12].sbox/U99  ( .A(\e/w[3][11] ), .B(\e/w[3][10] ), .Z(n3056)
         );
  XOR \e/a/SBOX[12].sbox/U98  ( .A(\e/w[3][13] ), .B(n3095), .Z(
        \e/a/SBOX[12].sbox/y[16] ) );
  XOR \e/a/SBOX[12].sbox/U97  ( .A(\e/a/SBOX[12].sbox/y[16] ), .B(n3057), .Z(
        n3096) );
  XOR \e/a/SBOX[12].sbox/U96  ( .A(\e/a/SBOX[12].sbox/t[12] ), .B(
        \e/a/SBOX[12].sbox/t[15] ), .Z(n3057) );
  XOR \e/a/SBOX[12].sbox/U95  ( .A(n3096), .B(n3058), .Z(
        \e/a/SBOX[12].sbox/t[29] ) );
  XOR \e/a/SBOX[12].sbox/U94  ( .A(\e/a/SBOX[12].sbox/t[28] ), .B(n3097), .Z(
        n3058) );
  XOR \e/a/SBOX[12].sbox/U93  ( .A(\e/w[3][8] ), .B(n3059), .Z(
        \e/a/SBOX[12].sbox/y[1] ) );
  XOR \e/a/SBOX[12].sbox/U92  ( .A(\e/w[3][14] ), .B(\e/w[3][13] ), .Z(n3059)
         );
  XOR \e/a/SBOX[12].sbox/U91  ( .A(\e/w[3][15] ), .B(\e/a/SBOX[12].sbox/y[1] ), 
        .Z(\e/a/SBOX[12].sbox/y[2] ) );
  XOR \e/a/SBOX[12].sbox/U90  ( .A(n3061), .B(n3060), .Z(
        \e/a/SBOX[12].sbox/t[25] ) );
  XOR \e/a/SBOX[12].sbox/U89  ( .A(n3063), .B(n3062), .Z(n3060) );
  XOR \e/a/SBOX[12].sbox/U88  ( .A(\e/w[3][15] ), .B(\e/w[3][13] ), .Z(n3061)
         );
  XOR \e/a/SBOX[12].sbox/U87  ( .A(\e/a/SBOX[12].sbox/t[13] ), .B(
        \e/a/SBOX[12].sbox/t[15] ), .Z(n3062) );
  XOR \e/a/SBOX[12].sbox/U86  ( .A(\e/a/SBOX[12].sbox/t[3] ), .B(
        \e/a/SBOX[12].sbox/t[5] ), .Z(n3063) );
  XOR \e/a/SBOX[12].sbox/U85  ( .A(\e/a/SBOX[12].sbox/t[39] ), .B(
        \e/a/SBOX[12].sbox/t[25] ), .Z(\e/a/SBOX[12].sbox/t[40] ) );
  XOR \e/a/SBOX[12].sbox/U84  ( .A(\e/w[3][9] ), .B(\e/a/SBOX[12].sbox/y[1] ), 
        .Z(\e/a/SBOX[12].sbox/y[5] ) );
  XOR \e/a/SBOX[12].sbox/U83  ( .A(n3065), .B(n3064), .Z(
        \e/a/SBOX[12].sbox/y[15] ) );
  XOR \e/a/SBOX[12].sbox/U82  ( .A(\e/w[3][11] ), .B(\e/w[3][9] ), .Z(n3064)
         );
  XOR \e/a/SBOX[12].sbox/U81  ( .A(\e/w[3][15] ), .B(\e/w[3][12] ), .Z(n3065)
         );
  XOR \e/a/SBOX[12].sbox/U80  ( .A(n3067), .B(n3066), .Z(
        \e/a/SBOX[12].sbox/t[21] ) );
  XOR \e/a/SBOX[12].sbox/U79  ( .A(n3069), .B(n3068), .Z(n3066) );
  XOR \e/a/SBOX[12].sbox/U78  ( .A(\e/a/SBOX[12].sbox/y[15] ), .B(n3092), .Z(
        n3067) );
  XOR \e/a/SBOX[12].sbox/U77  ( .A(\e/a/SBOX[12].sbox/t[13] ), .B(\e/w[3][10] ), .Z(n3068) );
  XOR \e/a/SBOX[12].sbox/U76  ( .A(\e/a/SBOX[12].sbox/t[3] ), .B(
        \e/a/SBOX[12].sbox/t[12] ), .Z(n3069) );
  XOR \e/a/SBOX[12].sbox/U75  ( .A(\e/a/SBOX[12].sbox/t[21] ), .B(n3070), .Z(
        \e/a/SBOX[12].sbox/t[43] ) );
  XOR \e/a/SBOX[12].sbox/U74  ( .A(\e/a/SBOX[12].sbox/t[28] ), .B(
        \e/a/SBOX[12].sbox/t[39] ), .Z(n3070) );
  XOR \e/a/SBOX[12].sbox/U73  ( .A(n3096), .B(n3093), .Z(
        \e/a/SBOX[12].sbox/t[24] ) );
  XOR \e/a/SBOX[12].sbox/U72  ( .A(\e/a/SBOX[12].sbox/t[32] ), .B(
        \e/a/SBOX[12].sbox/t[24] ), .Z(\e/a/SBOX[12].sbox/t[33] ) );
  XOR \e/a/SBOX[12].sbox/U71  ( .A(\e/w[3][12] ), .B(\e/a/SBOX[12].sbox/y[1] ), 
        .Z(\e/a/SBOX[12].sbox/y[4] ) );
  XOR \e/a/SBOX[12].sbox/U70  ( .A(n3072), .B(n3071), .Z(
        \e/a/SBOX[12].sbox/t[30] ) );
  XOR \e/a/SBOX[12].sbox/U69  ( .A(\e/w[3][9] ), .B(n3073), .Z(n3071) );
  XOR \e/a/SBOX[12].sbox/U68  ( .A(\e/a/SBOX[12].sbox/t[13] ), .B(
        \e/a/SBOX[12].sbox/t[15] ), .Z(n3072) );
  XOR \e/a/SBOX[12].sbox/U67  ( .A(\e/a/SBOX[12].sbox/t[8] ), .B(
        \e/a/SBOX[12].sbox/t[10] ), .Z(n3073) );
  XOR \e/a/SBOX[12].sbox/U66  ( .A(\e/a/SBOX[12].sbox/t[30] ), .B(n3074), .Z(
        \e/a/SBOX[12].sbox/t[37] ) );
  XOR \e/a/SBOX[12].sbox/U65  ( .A(\e/a/SBOX[12].sbox/t[32] ), .B(
        \e/a/SBOX[12].sbox/t[36] ), .Z(n3074) );
  XOR \e/a/SBOX[12].sbox/U64  ( .A(\e/w[3][15] ), .B(\e/w[3][10] ), .Z(n3094)
         );
  XOR \e/a/SBOX[12].sbox/U63  ( .A(\e/a/SBOX[12].sbox/y[5] ), .B(n3094), .Z(
        \e/a/SBOX[12].sbox/y[3] ) );
  XOR \e/a/SBOX[12].sbox/U62  ( .A(n3076), .B(n3075), .Z(
        \e/a/SBOX[12].sbox/t[23] ) );
  XOR \e/a/SBOX[12].sbox/U61  ( .A(n3078), .B(n3077), .Z(n3075) );
  XOR \e/a/SBOX[12].sbox/U60  ( .A(n3094), .B(n3079), .Z(n3076) );
  XOR \e/a/SBOX[12].sbox/U59  ( .A(\e/w[3][13] ), .B(\e/w[3][11] ), .Z(n3077)
         );
  XOR \e/a/SBOX[12].sbox/U58  ( .A(\e/a/SBOX[12].sbox/t[12] ), .B(
        \e/a/SBOX[12].sbox/t[13] ), .Z(n3078) );
  XOR \e/a/SBOX[12].sbox/U57  ( .A(\e/a/SBOX[12].sbox/t[7] ), .B(
        \e/a/SBOX[12].sbox/t[8] ), .Z(n3079) );
  XOR \e/a/SBOX[12].sbox/U56  ( .A(\e/a/SBOX[12].sbox/t[36] ), .B(
        \e/a/SBOX[12].sbox/t[23] ), .Z(\e/a/SBOX[12].sbox/t[44] ) );
  XOR \e/a/SBOX[12].sbox/U55  ( .A(n3094), .B(n3080), .Z(
        \e/a/SBOX[12].sbox/y[12] ) );
  XOR \e/a/SBOX[12].sbox/U54  ( .A(\e/w[3][12] ), .B(\e/w[3][9] ), .Z(n3080)
         );
  XOR \e/a/SBOX[12].sbox/U53  ( .A(\e/a/SBOX[12].sbox/y[15] ), .B(n3081), .Z(
        \e/a/SBOX[12].sbox/y[10] ) );
  XOR \e/a/SBOX[12].sbox/U52  ( .A(\e/w[3][14] ), .B(\e/w[3][13] ), .Z(n3081)
         );
  XOR \e/a/SBOX[12].sbox/U51  ( .A(n3094), .B(n3082), .Z(
        \e/a/SBOX[12].sbox/y[17] ) );
  XOR \e/a/SBOX[12].sbox/U50  ( .A(\e/w[3][13] ), .B(\e/w[3][12] ), .Z(n3082)
         );
  XOR \e/a/SBOX[12].sbox/U49  ( .A(\e/w[3][14] ), .B(n3095), .Z(
        \e/a/SBOX[12].sbox/y[11] ) );
  XOR \e/a/SBOX[12].sbox/U48  ( .A(\e/w[3][8] ), .B(\e/a/SBOX[12].sbox/y[11] ), 
        .Z(\e/a/SBOX[12].sbox/y[7] ) );
  XOR \e/a/SBOX[12].sbox/U47  ( .A(\e/w[3][8] ), .B(\e/a/SBOX[12].sbox/y[15] ), 
        .Z(\e/a/SBOX[12].sbox/y[6] ) );
  XOR \e/a/SBOX[12].sbox/U46  ( .A(\e/a/SBOX[12].sbox/t[26] ), .B(
        \e/a/SBOX[12].sbox/t[24] ), .Z(\e/a/SBOX[12].sbox/t[27] ) );
  XOR \e/a/SBOX[12].sbox/U45  ( .A(\e/a/SBOX[12].sbox/t[36] ), .B(
        \e/a/SBOX[12].sbox/t[27] ), .Z(\e/a/SBOX[12].sbox/t[38] ) );
  XOR \e/a/SBOX[12].sbox/U44  ( .A(n3096), .B(n3083), .Z(
        \e/a/SBOX[12].sbox/t[31] ) );
  XOR \e/a/SBOX[12].sbox/U43  ( .A(\e/a/SBOX[12].sbox/t[26] ), .B(n3097), .Z(
        n3083) );
  XOR \b/SBOX[15].sbox/U157  ( .A(\b/SBOX[15].sbox/z[12] ), .B(n2940), .Z(
        n3004) );
  XOR \b/SBOX[15].sbox/U156  ( .A(\b/SBOX[15].sbox/z[0] ), .B(
        \b/SBOX[15].sbox/z[2] ), .Z(n2940) );
  XOR \b/SBOX[15].sbox/U155  ( .A(n2942), .B(n2941), .Z(n3003) );
  XOR \b/SBOX[15].sbox/U154  ( .A(\b/SBOX[15].sbox/z[15] ), .B(
        \b/SBOX[15].sbox/z[16] ), .Z(n2941) );
  XOR \b/SBOX[15].sbox/U153  ( .A(\b/SBOX[15].sbox/z[5] ), .B(
        \b/SBOX[15].sbox/z[13] ), .Z(n2942) );
  XOR \b/SBOX[15].sbox/U152  ( .A(n3003), .B(n2943), .Z(n3017) );
  XOR \b/SBOX[15].sbox/U151  ( .A(\b/SBOX[15].sbox/z[3] ), .B(n3004), .Z(n2943) );
  XOR \b/SBOX[15].sbox/U150  ( .A(n2945), .B(n2944), .Z(n3018) );
  XOR \b/SBOX[15].sbox/U149  ( .A(n3003), .B(n2946), .Z(n2944) );
  XOR \b/SBOX[15].sbox/U148  ( .A(\b/SBOX[15].sbox/z[8] ), .B(
        \b/SBOX[15].sbox/z[12] ), .Z(n2945) );
  XOR \b/SBOX[15].sbox/U147  ( .A(\b/SBOX[15].sbox/z[4] ), .B(
        \b/SBOX[15].sbox/z[7] ), .Z(n2946) );
  XOR \b/SBOX[15].sbox/U146  ( .A(n3004), .B(n2947), .Z(n3006) );
  XOR \b/SBOX[15].sbox/U145  ( .A(\b/SBOX[15].sbox/z[8] ), .B(
        \b/SBOX[15].sbox/z[14] ), .Z(n2947) );
  XOR \b/SBOX[15].sbox/U144  ( .A(n2949), .B(n2948), .Z(n3019) );
  XOR \b/SBOX[15].sbox/U143  ( .A(\b/SBOX[15].sbox/z[17] ), .B(n3006), .Z(
        n2948) );
  XOR \b/SBOX[15].sbox/U142  ( .A(\b/SBOX[15].sbox/z[6] ), .B(
        \b/SBOX[15].sbox/z[15] ), .Z(n2949) );
  XOR \b/SBOX[15].sbox/U141  ( .A(\b/SBOX[15].sbox/z[9] ), .B(n2950), .Z(n3007) );
  XOR \b/SBOX[15].sbox/U140  ( .A(\b/SBOX[15].sbox/z[0] ), .B(
        \b/SBOX[15].sbox/z[1] ), .Z(n2950) );
  XOR \b/SBOX[15].sbox/U139  ( .A(\b/SBOX[15].sbox/z[16] ), .B(n2951), .Z(
        n3005) );
  XOR \b/SBOX[15].sbox/U138  ( .A(\b/SBOX[15].sbox/z[10] ), .B(
        \b/SBOX[15].sbox/z[15] ), .Z(n2951) );
  XOR \b/SBOX[15].sbox/U137  ( .A(n2953), .B(n2952), .Z(n3020) );
  XOR \b/SBOX[15].sbox/U136  ( .A(n3007), .B(n3005), .Z(n2952) );
  XOR \b/SBOX[15].sbox/U135  ( .A(\b/SBOX[15].sbox/z[6] ), .B(
        \b/SBOX[15].sbox/z[7] ), .Z(n2953) );
  XOR \b/SBOX[15].sbox/U134  ( .A(\b/SBOX[15].sbox/z[4] ), .B(n3005), .Z(n3008) );
  XOR \b/SBOX[15].sbox/U133  ( .A(n3008), .B(n2954), .Z(n3009) );
  XOR \b/SBOX[15].sbox/U132  ( .A(\b/SBOX[15].sbox/z[3] ), .B(
        \b/SBOX[15].sbox/z[7] ), .Z(n2954) );
  XOR \b/SBOX[15].sbox/U131  ( .A(n3006), .B(n2955), .Z(shift_row_out[26]) );
  XOR \b/SBOX[15].sbox/U130  ( .A(\b/SBOX[15].sbox/z[11] ), .B(n3009), .Z(
        n2955) );
  XOR \b/SBOX[15].sbox/U129  ( .A(n2957), .B(n2956), .Z(shift_row_out[27]) );
  XOR \b/SBOX[15].sbox/U128  ( .A(n3008), .B(n2958), .Z(n2956) );
  XOR \b/SBOX[15].sbox/U127  ( .A(\b/SBOX[15].sbox/z[5] ), .B(
        \b/SBOX[15].sbox/z[9] ), .Z(n2957) );
  XOR \b/SBOX[15].sbox/U126  ( .A(\b/SBOX[15].sbox/z[1] ), .B(
        \b/SBOX[15].sbox/z[2] ), .Z(n2958) );
  XOR \b/SBOX[15].sbox/U125  ( .A(n3007), .B(n2959), .Z(shift_row_out[28]) );
  XOR \b/SBOX[15].sbox/U124  ( .A(\b/SBOX[15].sbox/z[3] ), .B(n3008), .Z(n2959) );
  XOR \b/SBOX[15].sbox/U123  ( .A(n3009), .B(n2960), .Z(shift_row_out[31]) );
  XOR \b/SBOX[15].sbox/U122  ( .A(\b/SBOX[15].sbox/z[6] ), .B(
        \b/SBOX[15].sbox/z[9] ), .Z(n2960) );
  XOR \b/SBOX[15].sbox/U121  ( .A(n2962), .B(n2961), .Z(n3010) );
  XOR \b/SBOX[15].sbox/U120  ( .A(n2964), .B(n2963), .Z(n2961) );
  XOR \b/SBOX[15].sbox/U119  ( .A(msg[125]), .B(msg[121]), .Z(n2962) );
  XOR \b/SBOX[15].sbox/U118  ( .A(\b/SBOX[15].sbox/t[36] ), .B(
        \b/SBOX[15].sbox/t[39] ), .Z(n2963) );
  XOR \b/SBOX[15].sbox/U117  ( .A(\b/SBOX[15].sbox/t[3] ), .B(
        \b/SBOX[15].sbox/t[8] ), .Z(n2964) );
  XOR \b/SBOX[15].sbox/U116  ( .A(n2966), .B(n2965), .Z(
        \b/SBOX[15].sbox/t[41] ) );
  XOR \b/SBOX[15].sbox/U115  ( .A(n3010), .B(n2967), .Z(n2965) );
  XOR \b/SBOX[15].sbox/U114  ( .A(\b/SBOX[15].sbox/t[32] ), .B(msg[127]), .Z(
        n2966) );
  XOR \b/SBOX[15].sbox/U113  ( .A(\b/SBOX[15].sbox/t[5] ), .B(
        \b/SBOX[15].sbox/t[10] ), .Z(n2967) );
  XOR \b/SBOX[15].sbox/U112  ( .A(\b/SBOX[15].sbox/t[2] ), .B(msg[126]), .Z(
        n3011) );
  XOR \b/SBOX[15].sbox/U111  ( .A(n2969), .B(n2968), .Z(
        \b/SBOX[15].sbox/t[45] ) );
  XOR \b/SBOX[15].sbox/U110  ( .A(n3011), .B(n2970), .Z(n2968) );
  XOR \b/SBOX[15].sbox/U109  ( .A(msg[124]), .B(n3010), .Z(n2969) );
  XOR \b/SBOX[15].sbox/U108  ( .A(\b/SBOX[15].sbox/t[7] ), .B(
        \b/SBOX[15].sbox/t[28] ), .Z(n2970) );
  XOR \b/SBOX[15].sbox/U107  ( .A(n3011), .B(n2971), .Z(n3016) );
  XOR \b/SBOX[15].sbox/U106  ( .A(\b/SBOX[15].sbox/t[5] ), .B(msg[124]), .Z(
        n2971) );
  XOR \b/SBOX[15].sbox/U105  ( .A(msg[127]), .B(n2972), .Z(n3012) );
  XOR \b/SBOX[15].sbox/U104  ( .A(\b/SBOX[15].sbox/t[7] ), .B(
        \b/SBOX[15].sbox/t[10] ), .Z(n2972) );
  XOR \b/SBOX[15].sbox/U103  ( .A(n2974), .B(n2973), .Z(
        \b/SBOX[15].sbox/t[42] ) );
  XOR \b/SBOX[15].sbox/U102  ( .A(n3016), .B(n3012), .Z(n2973) );
  XOR \b/SBOX[15].sbox/U101  ( .A(\b/SBOX[15].sbox/t[28] ), .B(
        \b/SBOX[15].sbox/t[32] ), .Z(n2974) );
  XOR \b/SBOX[15].sbox/U100  ( .A(msg[121]), .B(n2975), .Z(n3014) );
  XOR \b/SBOX[15].sbox/U99  ( .A(msg[123]), .B(msg[122]), .Z(n2975) );
  XOR \b/SBOX[15].sbox/U98  ( .A(msg[125]), .B(n3014), .Z(
        \b/SBOX[15].sbox/y[16] ) );
  XOR \b/SBOX[15].sbox/U97  ( .A(\b/SBOX[15].sbox/y[16] ), .B(n2976), .Z(n3015) );
  XOR \b/SBOX[15].sbox/U96  ( .A(\b/SBOX[15].sbox/t[12] ), .B(
        \b/SBOX[15].sbox/t[15] ), .Z(n2976) );
  XOR \b/SBOX[15].sbox/U95  ( .A(n3015), .B(n2977), .Z(\b/SBOX[15].sbox/t[29] ) );
  XOR \b/SBOX[15].sbox/U94  ( .A(\b/SBOX[15].sbox/t[28] ), .B(n3016), .Z(n2977) );
  XOR \b/SBOX[15].sbox/U93  ( .A(msg[120]), .B(n2978), .Z(
        \b/SBOX[15].sbox/y[1] ) );
  XOR \b/SBOX[15].sbox/U92  ( .A(msg[126]), .B(msg[125]), .Z(n2978) );
  XOR \b/SBOX[15].sbox/U91  ( .A(msg[127]), .B(\b/SBOX[15].sbox/y[1] ), .Z(
        \b/SBOX[15].sbox/y[2] ) );
  XOR \b/SBOX[15].sbox/U90  ( .A(n2980), .B(n2979), .Z(\b/SBOX[15].sbox/t[25] ) );
  XOR \b/SBOX[15].sbox/U89  ( .A(n2982), .B(n2981), .Z(n2979) );
  XOR \b/SBOX[15].sbox/U88  ( .A(msg[127]), .B(msg[125]), .Z(n2980) );
  XOR \b/SBOX[15].sbox/U87  ( .A(\b/SBOX[15].sbox/t[13] ), .B(
        \b/SBOX[15].sbox/t[15] ), .Z(n2981) );
  XOR \b/SBOX[15].sbox/U86  ( .A(\b/SBOX[15].sbox/t[3] ), .B(
        \b/SBOX[15].sbox/t[5] ), .Z(n2982) );
  XOR \b/SBOX[15].sbox/U85  ( .A(\b/SBOX[15].sbox/t[39] ), .B(
        \b/SBOX[15].sbox/t[25] ), .Z(\b/SBOX[15].sbox/t[40] ) );
  XOR \b/SBOX[15].sbox/U84  ( .A(msg[121]), .B(\b/SBOX[15].sbox/y[1] ), .Z(
        \b/SBOX[15].sbox/y[5] ) );
  XOR \b/SBOX[15].sbox/U83  ( .A(n2984), .B(n2983), .Z(\b/SBOX[15].sbox/y[15] ) );
  XOR \b/SBOX[15].sbox/U82  ( .A(msg[123]), .B(msg[121]), .Z(n2983) );
  XOR \b/SBOX[15].sbox/U81  ( .A(msg[127]), .B(msg[124]), .Z(n2984) );
  XOR \b/SBOX[15].sbox/U80  ( .A(n2986), .B(n2985), .Z(\b/SBOX[15].sbox/t[21] ) );
  XOR \b/SBOX[15].sbox/U79  ( .A(n2988), .B(n2987), .Z(n2985) );
  XOR \b/SBOX[15].sbox/U78  ( .A(\b/SBOX[15].sbox/y[15] ), .B(n3011), .Z(n2986) );
  XOR \b/SBOX[15].sbox/U77  ( .A(\b/SBOX[15].sbox/t[13] ), .B(msg[122]), .Z(
        n2987) );
  XOR \b/SBOX[15].sbox/U76  ( .A(\b/SBOX[15].sbox/t[3] ), .B(
        \b/SBOX[15].sbox/t[12] ), .Z(n2988) );
  XOR \b/SBOX[15].sbox/U75  ( .A(\b/SBOX[15].sbox/t[21] ), .B(n2989), .Z(
        \b/SBOX[15].sbox/t[43] ) );
  XOR \b/SBOX[15].sbox/U74  ( .A(\b/SBOX[15].sbox/t[28] ), .B(
        \b/SBOX[15].sbox/t[39] ), .Z(n2989) );
  XOR \b/SBOX[15].sbox/U73  ( .A(n3015), .B(n3012), .Z(\b/SBOX[15].sbox/t[24] ) );
  XOR \b/SBOX[15].sbox/U72  ( .A(\b/SBOX[15].sbox/t[32] ), .B(
        \b/SBOX[15].sbox/t[24] ), .Z(\b/SBOX[15].sbox/t[33] ) );
  XOR \b/SBOX[15].sbox/U71  ( .A(msg[124]), .B(\b/SBOX[15].sbox/y[1] ), .Z(
        \b/SBOX[15].sbox/y[4] ) );
  XOR \b/SBOX[15].sbox/U70  ( .A(n2991), .B(n2990), .Z(\b/SBOX[15].sbox/t[30] ) );
  XOR \b/SBOX[15].sbox/U69  ( .A(msg[121]), .B(n2992), .Z(n2990) );
  XOR \b/SBOX[15].sbox/U68  ( .A(\b/SBOX[15].sbox/t[13] ), .B(
        \b/SBOX[15].sbox/t[15] ), .Z(n2991) );
  XOR \b/SBOX[15].sbox/U67  ( .A(\b/SBOX[15].sbox/t[8] ), .B(
        \b/SBOX[15].sbox/t[10] ), .Z(n2992) );
  XOR \b/SBOX[15].sbox/U66  ( .A(\b/SBOX[15].sbox/t[30] ), .B(n2993), .Z(
        \b/SBOX[15].sbox/t[37] ) );
  XOR \b/SBOX[15].sbox/U65  ( .A(\b/SBOX[15].sbox/t[32] ), .B(
        \b/SBOX[15].sbox/t[36] ), .Z(n2993) );
  XOR \b/SBOX[15].sbox/U64  ( .A(msg[127]), .B(msg[122]), .Z(n3013) );
  XOR \b/SBOX[15].sbox/U63  ( .A(\b/SBOX[15].sbox/y[5] ), .B(n3013), .Z(
        \b/SBOX[15].sbox/y[3] ) );
  XOR \b/SBOX[15].sbox/U62  ( .A(n2995), .B(n2994), .Z(\b/SBOX[15].sbox/t[23] ) );
  XOR \b/SBOX[15].sbox/U61  ( .A(n2997), .B(n2996), .Z(n2994) );
  XOR \b/SBOX[15].sbox/U60  ( .A(n3013), .B(n2998), .Z(n2995) );
  XOR \b/SBOX[15].sbox/U59  ( .A(msg[125]), .B(msg[123]), .Z(n2996) );
  XOR \b/SBOX[15].sbox/U58  ( .A(\b/SBOX[15].sbox/t[12] ), .B(
        \b/SBOX[15].sbox/t[13] ), .Z(n2997) );
  XOR \b/SBOX[15].sbox/U57  ( .A(\b/SBOX[15].sbox/t[7] ), .B(
        \b/SBOX[15].sbox/t[8] ), .Z(n2998) );
  XOR \b/SBOX[15].sbox/U56  ( .A(\b/SBOX[15].sbox/t[36] ), .B(
        \b/SBOX[15].sbox/t[23] ), .Z(\b/SBOX[15].sbox/t[44] ) );
  XOR \b/SBOX[15].sbox/U55  ( .A(n3013), .B(n2999), .Z(\b/SBOX[15].sbox/y[12] ) );
  XOR \b/SBOX[15].sbox/U54  ( .A(msg[124]), .B(msg[121]), .Z(n2999) );
  XOR \b/SBOX[15].sbox/U53  ( .A(\b/SBOX[15].sbox/y[15] ), .B(n3000), .Z(
        \b/SBOX[15].sbox/y[10] ) );
  XOR \b/SBOX[15].sbox/U52  ( .A(msg[126]), .B(msg[125]), .Z(n3000) );
  XOR \b/SBOX[15].sbox/U51  ( .A(n3013), .B(n3001), .Z(\b/SBOX[15].sbox/y[17] ) );
  XOR \b/SBOX[15].sbox/U50  ( .A(msg[125]), .B(msg[124]), .Z(n3001) );
  XOR \b/SBOX[15].sbox/U49  ( .A(msg[126]), .B(n3014), .Z(
        \b/SBOX[15].sbox/y[11] ) );
  XOR \b/SBOX[15].sbox/U48  ( .A(msg[120]), .B(\b/SBOX[15].sbox/y[11] ), .Z(
        \b/SBOX[15].sbox/y[7] ) );
  XOR \b/SBOX[15].sbox/U47  ( .A(msg[120]), .B(\b/SBOX[15].sbox/y[15] ), .Z(
        \b/SBOX[15].sbox/y[6] ) );
  XOR \b/SBOX[15].sbox/U46  ( .A(\b/SBOX[15].sbox/t[26] ), .B(
        \b/SBOX[15].sbox/t[24] ), .Z(\b/SBOX[15].sbox/t[27] ) );
  XOR \b/SBOX[15].sbox/U45  ( .A(\b/SBOX[15].sbox/t[36] ), .B(
        \b/SBOX[15].sbox/t[27] ), .Z(\b/SBOX[15].sbox/t[38] ) );
  XOR \b/SBOX[15].sbox/U44  ( .A(n3015), .B(n3002), .Z(\b/SBOX[15].sbox/t[31] ) );
  XOR \b/SBOX[15].sbox/U43  ( .A(\b/SBOX[15].sbox/t[26] ), .B(n3016), .Z(n3002) );
  XOR \b/SBOX[14].sbox/U157  ( .A(\b/SBOX[14].sbox/z[12] ), .B(n2859), .Z(
        n2923) );
  XOR \b/SBOX[14].sbox/U156  ( .A(\b/SBOX[14].sbox/z[0] ), .B(
        \b/SBOX[14].sbox/z[2] ), .Z(n2859) );
  XOR \b/SBOX[14].sbox/U155  ( .A(n2861), .B(n2860), .Z(n2922) );
  XOR \b/SBOX[14].sbox/U154  ( .A(\b/SBOX[14].sbox/z[15] ), .B(
        \b/SBOX[14].sbox/z[16] ), .Z(n2860) );
  XOR \b/SBOX[14].sbox/U153  ( .A(\b/SBOX[14].sbox/z[5] ), .B(
        \b/SBOX[14].sbox/z[13] ), .Z(n2861) );
  XOR \b/SBOX[14].sbox/U152  ( .A(n2922), .B(n2862), .Z(n2936) );
  XOR \b/SBOX[14].sbox/U151  ( .A(\b/SBOX[14].sbox/z[3] ), .B(n2923), .Z(n2862) );
  XOR \b/SBOX[14].sbox/U150  ( .A(n2864), .B(n2863), .Z(n2937) );
  XOR \b/SBOX[14].sbox/U149  ( .A(n2922), .B(n2865), .Z(n2863) );
  XOR \b/SBOX[14].sbox/U148  ( .A(\b/SBOX[14].sbox/z[8] ), .B(
        \b/SBOX[14].sbox/z[12] ), .Z(n2864) );
  XOR \b/SBOX[14].sbox/U147  ( .A(\b/SBOX[14].sbox/z[4] ), .B(
        \b/SBOX[14].sbox/z[7] ), .Z(n2865) );
  XOR \b/SBOX[14].sbox/U146  ( .A(n2923), .B(n2866), .Z(n2925) );
  XOR \b/SBOX[14].sbox/U145  ( .A(\b/SBOX[14].sbox/z[8] ), .B(
        \b/SBOX[14].sbox/z[14] ), .Z(n2866) );
  XOR \b/SBOX[14].sbox/U144  ( .A(n2868), .B(n2867), .Z(n2938) );
  XOR \b/SBOX[14].sbox/U143  ( .A(\b/SBOX[14].sbox/z[17] ), .B(n2925), .Z(
        n2867) );
  XOR \b/SBOX[14].sbox/U142  ( .A(\b/SBOX[14].sbox/z[6] ), .B(
        \b/SBOX[14].sbox/z[15] ), .Z(n2868) );
  XOR \b/SBOX[14].sbox/U141  ( .A(\b/SBOX[14].sbox/z[9] ), .B(n2869), .Z(n2926) );
  XOR \b/SBOX[14].sbox/U140  ( .A(\b/SBOX[14].sbox/z[0] ), .B(
        \b/SBOX[14].sbox/z[1] ), .Z(n2869) );
  XOR \b/SBOX[14].sbox/U139  ( .A(\b/SBOX[14].sbox/z[16] ), .B(n2870), .Z(
        n2924) );
  XOR \b/SBOX[14].sbox/U138  ( .A(\b/SBOX[14].sbox/z[10] ), .B(
        \b/SBOX[14].sbox/z[15] ), .Z(n2870) );
  XOR \b/SBOX[14].sbox/U137  ( .A(n2872), .B(n2871), .Z(n2939) );
  XOR \b/SBOX[14].sbox/U136  ( .A(n2926), .B(n2924), .Z(n2871) );
  XOR \b/SBOX[14].sbox/U135  ( .A(\b/SBOX[14].sbox/z[6] ), .B(
        \b/SBOX[14].sbox/z[7] ), .Z(n2872) );
  XOR \b/SBOX[14].sbox/U134  ( .A(\b/SBOX[14].sbox/z[4] ), .B(n2924), .Z(n2927) );
  XOR \b/SBOX[14].sbox/U133  ( .A(n2927), .B(n2873), .Z(n2928) );
  XOR \b/SBOX[14].sbox/U132  ( .A(\b/SBOX[14].sbox/z[3] ), .B(
        \b/SBOX[14].sbox/z[7] ), .Z(n2873) );
  XOR \b/SBOX[14].sbox/U131  ( .A(n2925), .B(n2874), .Z(shift_row_out[50]) );
  XOR \b/SBOX[14].sbox/U130  ( .A(\b/SBOX[14].sbox/z[11] ), .B(n2928), .Z(
        n2874) );
  XOR \b/SBOX[14].sbox/U129  ( .A(n2876), .B(n2875), .Z(shift_row_out[51]) );
  XOR \b/SBOX[14].sbox/U128  ( .A(n2927), .B(n2877), .Z(n2875) );
  XOR \b/SBOX[14].sbox/U127  ( .A(\b/SBOX[14].sbox/z[5] ), .B(
        \b/SBOX[14].sbox/z[9] ), .Z(n2876) );
  XOR \b/SBOX[14].sbox/U126  ( .A(\b/SBOX[14].sbox/z[1] ), .B(
        \b/SBOX[14].sbox/z[2] ), .Z(n2877) );
  XOR \b/SBOX[14].sbox/U125  ( .A(n2926), .B(n2878), .Z(shift_row_out[52]) );
  XOR \b/SBOX[14].sbox/U124  ( .A(\b/SBOX[14].sbox/z[3] ), .B(n2927), .Z(n2878) );
  XOR \b/SBOX[14].sbox/U123  ( .A(n2928), .B(n2879), .Z(shift_row_out[55]) );
  XOR \b/SBOX[14].sbox/U122  ( .A(\b/SBOX[14].sbox/z[6] ), .B(
        \b/SBOX[14].sbox/z[9] ), .Z(n2879) );
  XOR \b/SBOX[14].sbox/U121  ( .A(n2881), .B(n2880), .Z(n2929) );
  XOR \b/SBOX[14].sbox/U120  ( .A(n2883), .B(n2882), .Z(n2880) );
  XOR \b/SBOX[14].sbox/U119  ( .A(msg[117]), .B(msg[113]), .Z(n2881) );
  XOR \b/SBOX[14].sbox/U118  ( .A(\b/SBOX[14].sbox/t[36] ), .B(
        \b/SBOX[14].sbox/t[39] ), .Z(n2882) );
  XOR \b/SBOX[14].sbox/U117  ( .A(\b/SBOX[14].sbox/t[3] ), .B(
        \b/SBOX[14].sbox/t[8] ), .Z(n2883) );
  XOR \b/SBOX[14].sbox/U116  ( .A(n2885), .B(n2884), .Z(
        \b/SBOX[14].sbox/t[41] ) );
  XOR \b/SBOX[14].sbox/U115  ( .A(n2929), .B(n2886), .Z(n2884) );
  XOR \b/SBOX[14].sbox/U114  ( .A(\b/SBOX[14].sbox/t[32] ), .B(msg[119]), .Z(
        n2885) );
  XOR \b/SBOX[14].sbox/U113  ( .A(\b/SBOX[14].sbox/t[5] ), .B(
        \b/SBOX[14].sbox/t[10] ), .Z(n2886) );
  XOR \b/SBOX[14].sbox/U112  ( .A(\b/SBOX[14].sbox/t[2] ), .B(msg[118]), .Z(
        n2930) );
  XOR \b/SBOX[14].sbox/U111  ( .A(n2888), .B(n2887), .Z(
        \b/SBOX[14].sbox/t[45] ) );
  XOR \b/SBOX[14].sbox/U110  ( .A(n2930), .B(n2889), .Z(n2887) );
  XOR \b/SBOX[14].sbox/U109  ( .A(msg[116]), .B(n2929), .Z(n2888) );
  XOR \b/SBOX[14].sbox/U108  ( .A(\b/SBOX[14].sbox/t[7] ), .B(
        \b/SBOX[14].sbox/t[28] ), .Z(n2889) );
  XOR \b/SBOX[14].sbox/U107  ( .A(n2930), .B(n2890), .Z(n2935) );
  XOR \b/SBOX[14].sbox/U106  ( .A(\b/SBOX[14].sbox/t[5] ), .B(msg[116]), .Z(
        n2890) );
  XOR \b/SBOX[14].sbox/U105  ( .A(msg[119]), .B(n2891), .Z(n2931) );
  XOR \b/SBOX[14].sbox/U104  ( .A(\b/SBOX[14].sbox/t[7] ), .B(
        \b/SBOX[14].sbox/t[10] ), .Z(n2891) );
  XOR \b/SBOX[14].sbox/U103  ( .A(n2893), .B(n2892), .Z(
        \b/SBOX[14].sbox/t[42] ) );
  XOR \b/SBOX[14].sbox/U102  ( .A(n2935), .B(n2931), .Z(n2892) );
  XOR \b/SBOX[14].sbox/U101  ( .A(\b/SBOX[14].sbox/t[28] ), .B(
        \b/SBOX[14].sbox/t[32] ), .Z(n2893) );
  XOR \b/SBOX[14].sbox/U100  ( .A(msg[113]), .B(n2894), .Z(n2933) );
  XOR \b/SBOX[14].sbox/U99  ( .A(msg[115]), .B(msg[114]), .Z(n2894) );
  XOR \b/SBOX[14].sbox/U98  ( .A(msg[117]), .B(n2933), .Z(
        \b/SBOX[14].sbox/y[16] ) );
  XOR \b/SBOX[14].sbox/U97  ( .A(\b/SBOX[14].sbox/y[16] ), .B(n2895), .Z(n2934) );
  XOR \b/SBOX[14].sbox/U96  ( .A(\b/SBOX[14].sbox/t[12] ), .B(
        \b/SBOX[14].sbox/t[15] ), .Z(n2895) );
  XOR \b/SBOX[14].sbox/U95  ( .A(n2934), .B(n2896), .Z(\b/SBOX[14].sbox/t[29] ) );
  XOR \b/SBOX[14].sbox/U94  ( .A(\b/SBOX[14].sbox/t[28] ), .B(n2935), .Z(n2896) );
  XOR \b/SBOX[14].sbox/U93  ( .A(msg[112]), .B(n2897), .Z(
        \b/SBOX[14].sbox/y[1] ) );
  XOR \b/SBOX[14].sbox/U92  ( .A(msg[118]), .B(msg[117]), .Z(n2897) );
  XOR \b/SBOX[14].sbox/U91  ( .A(msg[119]), .B(\b/SBOX[14].sbox/y[1] ), .Z(
        \b/SBOX[14].sbox/y[2] ) );
  XOR \b/SBOX[14].sbox/U90  ( .A(n2899), .B(n2898), .Z(\b/SBOX[14].sbox/t[25] ) );
  XOR \b/SBOX[14].sbox/U89  ( .A(n2901), .B(n2900), .Z(n2898) );
  XOR \b/SBOX[14].sbox/U88  ( .A(msg[119]), .B(msg[117]), .Z(n2899) );
  XOR \b/SBOX[14].sbox/U87  ( .A(\b/SBOX[14].sbox/t[13] ), .B(
        \b/SBOX[14].sbox/t[15] ), .Z(n2900) );
  XOR \b/SBOX[14].sbox/U86  ( .A(\b/SBOX[14].sbox/t[3] ), .B(
        \b/SBOX[14].sbox/t[5] ), .Z(n2901) );
  XOR \b/SBOX[14].sbox/U85  ( .A(\b/SBOX[14].sbox/t[39] ), .B(
        \b/SBOX[14].sbox/t[25] ), .Z(\b/SBOX[14].sbox/t[40] ) );
  XOR \b/SBOX[14].sbox/U84  ( .A(msg[113]), .B(\b/SBOX[14].sbox/y[1] ), .Z(
        \b/SBOX[14].sbox/y[5] ) );
  XOR \b/SBOX[14].sbox/U83  ( .A(n2903), .B(n2902), .Z(\b/SBOX[14].sbox/y[15] ) );
  XOR \b/SBOX[14].sbox/U82  ( .A(msg[115]), .B(msg[113]), .Z(n2902) );
  XOR \b/SBOX[14].sbox/U81  ( .A(msg[119]), .B(msg[116]), .Z(n2903) );
  XOR \b/SBOX[14].sbox/U80  ( .A(n2905), .B(n2904), .Z(\b/SBOX[14].sbox/t[21] ) );
  XOR \b/SBOX[14].sbox/U79  ( .A(n2907), .B(n2906), .Z(n2904) );
  XOR \b/SBOX[14].sbox/U78  ( .A(\b/SBOX[14].sbox/y[15] ), .B(n2930), .Z(n2905) );
  XOR \b/SBOX[14].sbox/U77  ( .A(\b/SBOX[14].sbox/t[13] ), .B(msg[114]), .Z(
        n2906) );
  XOR \b/SBOX[14].sbox/U76  ( .A(\b/SBOX[14].sbox/t[3] ), .B(
        \b/SBOX[14].sbox/t[12] ), .Z(n2907) );
  XOR \b/SBOX[14].sbox/U75  ( .A(\b/SBOX[14].sbox/t[21] ), .B(n2908), .Z(
        \b/SBOX[14].sbox/t[43] ) );
  XOR \b/SBOX[14].sbox/U74  ( .A(\b/SBOX[14].sbox/t[28] ), .B(
        \b/SBOX[14].sbox/t[39] ), .Z(n2908) );
  XOR \b/SBOX[14].sbox/U73  ( .A(n2934), .B(n2931), .Z(\b/SBOX[14].sbox/t[24] ) );
  XOR \b/SBOX[14].sbox/U72  ( .A(\b/SBOX[14].sbox/t[32] ), .B(
        \b/SBOX[14].sbox/t[24] ), .Z(\b/SBOX[14].sbox/t[33] ) );
  XOR \b/SBOX[14].sbox/U71  ( .A(msg[116]), .B(\b/SBOX[14].sbox/y[1] ), .Z(
        \b/SBOX[14].sbox/y[4] ) );
  XOR \b/SBOX[14].sbox/U70  ( .A(n2910), .B(n2909), .Z(\b/SBOX[14].sbox/t[30] ) );
  XOR \b/SBOX[14].sbox/U69  ( .A(msg[113]), .B(n2911), .Z(n2909) );
  XOR \b/SBOX[14].sbox/U68  ( .A(\b/SBOX[14].sbox/t[13] ), .B(
        \b/SBOX[14].sbox/t[15] ), .Z(n2910) );
  XOR \b/SBOX[14].sbox/U67  ( .A(\b/SBOX[14].sbox/t[8] ), .B(
        \b/SBOX[14].sbox/t[10] ), .Z(n2911) );
  XOR \b/SBOX[14].sbox/U66  ( .A(\b/SBOX[14].sbox/t[30] ), .B(n2912), .Z(
        \b/SBOX[14].sbox/t[37] ) );
  XOR \b/SBOX[14].sbox/U65  ( .A(\b/SBOX[14].sbox/t[32] ), .B(
        \b/SBOX[14].sbox/t[36] ), .Z(n2912) );
  XOR \b/SBOX[14].sbox/U64  ( .A(msg[119]), .B(msg[114]), .Z(n2932) );
  XOR \b/SBOX[14].sbox/U63  ( .A(\b/SBOX[14].sbox/y[5] ), .B(n2932), .Z(
        \b/SBOX[14].sbox/y[3] ) );
  XOR \b/SBOX[14].sbox/U62  ( .A(n2914), .B(n2913), .Z(\b/SBOX[14].sbox/t[23] ) );
  XOR \b/SBOX[14].sbox/U61  ( .A(n2916), .B(n2915), .Z(n2913) );
  XOR \b/SBOX[14].sbox/U60  ( .A(n2932), .B(n2917), .Z(n2914) );
  XOR \b/SBOX[14].sbox/U59  ( .A(msg[117]), .B(msg[115]), .Z(n2915) );
  XOR \b/SBOX[14].sbox/U58  ( .A(\b/SBOX[14].sbox/t[12] ), .B(
        \b/SBOX[14].sbox/t[13] ), .Z(n2916) );
  XOR \b/SBOX[14].sbox/U57  ( .A(\b/SBOX[14].sbox/t[7] ), .B(
        \b/SBOX[14].sbox/t[8] ), .Z(n2917) );
  XOR \b/SBOX[14].sbox/U56  ( .A(\b/SBOX[14].sbox/t[36] ), .B(
        \b/SBOX[14].sbox/t[23] ), .Z(\b/SBOX[14].sbox/t[44] ) );
  XOR \b/SBOX[14].sbox/U55  ( .A(n2932), .B(n2918), .Z(\b/SBOX[14].sbox/y[12] ) );
  XOR \b/SBOX[14].sbox/U54  ( .A(msg[116]), .B(msg[113]), .Z(n2918) );
  XOR \b/SBOX[14].sbox/U53  ( .A(\b/SBOX[14].sbox/y[15] ), .B(n2919), .Z(
        \b/SBOX[14].sbox/y[10] ) );
  XOR \b/SBOX[14].sbox/U52  ( .A(msg[118]), .B(msg[117]), .Z(n2919) );
  XOR \b/SBOX[14].sbox/U51  ( .A(n2932), .B(n2920), .Z(\b/SBOX[14].sbox/y[17] ) );
  XOR \b/SBOX[14].sbox/U50  ( .A(msg[117]), .B(msg[116]), .Z(n2920) );
  XOR \b/SBOX[14].sbox/U49  ( .A(msg[118]), .B(n2933), .Z(
        \b/SBOX[14].sbox/y[11] ) );
  XOR \b/SBOX[14].sbox/U48  ( .A(msg[112]), .B(\b/SBOX[14].sbox/y[11] ), .Z(
        \b/SBOX[14].sbox/y[7] ) );
  XOR \b/SBOX[14].sbox/U47  ( .A(msg[112]), .B(\b/SBOX[14].sbox/y[15] ), .Z(
        \b/SBOX[14].sbox/y[6] ) );
  XOR \b/SBOX[14].sbox/U46  ( .A(\b/SBOX[14].sbox/t[26] ), .B(
        \b/SBOX[14].sbox/t[24] ), .Z(\b/SBOX[14].sbox/t[27] ) );
  XOR \b/SBOX[14].sbox/U45  ( .A(\b/SBOX[14].sbox/t[36] ), .B(
        \b/SBOX[14].sbox/t[27] ), .Z(\b/SBOX[14].sbox/t[38] ) );
  XOR \b/SBOX[14].sbox/U44  ( .A(n2934), .B(n2921), .Z(\b/SBOX[14].sbox/t[31] ) );
  XOR \b/SBOX[14].sbox/U43  ( .A(\b/SBOX[14].sbox/t[26] ), .B(n2935), .Z(n2921) );
  XOR \b/SBOX[13].sbox/U157  ( .A(\b/SBOX[13].sbox/z[12] ), .B(n2778), .Z(
        n2842) );
  XOR \b/SBOX[13].sbox/U156  ( .A(\b/SBOX[13].sbox/z[0] ), .B(
        \b/SBOX[13].sbox/z[2] ), .Z(n2778) );
  XOR \b/SBOX[13].sbox/U155  ( .A(n2780), .B(n2779), .Z(n2841) );
  XOR \b/SBOX[13].sbox/U154  ( .A(\b/SBOX[13].sbox/z[15] ), .B(
        \b/SBOX[13].sbox/z[16] ), .Z(n2779) );
  XOR \b/SBOX[13].sbox/U153  ( .A(\b/SBOX[13].sbox/z[5] ), .B(
        \b/SBOX[13].sbox/z[13] ), .Z(n2780) );
  XOR \b/SBOX[13].sbox/U152  ( .A(n2841), .B(n2781), .Z(n2855) );
  XOR \b/SBOX[13].sbox/U151  ( .A(\b/SBOX[13].sbox/z[3] ), .B(n2842), .Z(n2781) );
  XOR \b/SBOX[13].sbox/U150  ( .A(n2783), .B(n2782), .Z(n2856) );
  XOR \b/SBOX[13].sbox/U149  ( .A(n2841), .B(n2784), .Z(n2782) );
  XOR \b/SBOX[13].sbox/U148  ( .A(\b/SBOX[13].sbox/z[8] ), .B(
        \b/SBOX[13].sbox/z[12] ), .Z(n2783) );
  XOR \b/SBOX[13].sbox/U147  ( .A(\b/SBOX[13].sbox/z[4] ), .B(
        \b/SBOX[13].sbox/z[7] ), .Z(n2784) );
  XOR \b/SBOX[13].sbox/U146  ( .A(n2842), .B(n2785), .Z(n2844) );
  XOR \b/SBOX[13].sbox/U145  ( .A(\b/SBOX[13].sbox/z[8] ), .B(
        \b/SBOX[13].sbox/z[14] ), .Z(n2785) );
  XOR \b/SBOX[13].sbox/U144  ( .A(n2787), .B(n2786), .Z(n2857) );
  XOR \b/SBOX[13].sbox/U143  ( .A(\b/SBOX[13].sbox/z[17] ), .B(n2844), .Z(
        n2786) );
  XOR \b/SBOX[13].sbox/U142  ( .A(\b/SBOX[13].sbox/z[6] ), .B(
        \b/SBOX[13].sbox/z[15] ), .Z(n2787) );
  XOR \b/SBOX[13].sbox/U141  ( .A(\b/SBOX[13].sbox/z[9] ), .B(n2788), .Z(n2845) );
  XOR \b/SBOX[13].sbox/U140  ( .A(\b/SBOX[13].sbox/z[0] ), .B(
        \b/SBOX[13].sbox/z[1] ), .Z(n2788) );
  XOR \b/SBOX[13].sbox/U139  ( .A(\b/SBOX[13].sbox/z[16] ), .B(n2789), .Z(
        n2843) );
  XOR \b/SBOX[13].sbox/U138  ( .A(\b/SBOX[13].sbox/z[10] ), .B(
        \b/SBOX[13].sbox/z[15] ), .Z(n2789) );
  XOR \b/SBOX[13].sbox/U137  ( .A(n2791), .B(n2790), .Z(n2858) );
  XOR \b/SBOX[13].sbox/U136  ( .A(n2845), .B(n2843), .Z(n2790) );
  XOR \b/SBOX[13].sbox/U135  ( .A(\b/SBOX[13].sbox/z[6] ), .B(
        \b/SBOX[13].sbox/z[7] ), .Z(n2791) );
  XOR \b/SBOX[13].sbox/U134  ( .A(\b/SBOX[13].sbox/z[4] ), .B(n2843), .Z(n2846) );
  XOR \b/SBOX[13].sbox/U133  ( .A(n2846), .B(n2792), .Z(n2847) );
  XOR \b/SBOX[13].sbox/U132  ( .A(\b/SBOX[13].sbox/z[3] ), .B(
        \b/SBOX[13].sbox/z[7] ), .Z(n2792) );
  XOR \b/SBOX[13].sbox/U131  ( .A(n2844), .B(n2793), .Z(shift_row_out[74]) );
  XOR \b/SBOX[13].sbox/U130  ( .A(\b/SBOX[13].sbox/z[11] ), .B(n2847), .Z(
        n2793) );
  XOR \b/SBOX[13].sbox/U129  ( .A(n2795), .B(n2794), .Z(shift_row_out[75]) );
  XOR \b/SBOX[13].sbox/U128  ( .A(n2846), .B(n2796), .Z(n2794) );
  XOR \b/SBOX[13].sbox/U127  ( .A(\b/SBOX[13].sbox/z[5] ), .B(
        \b/SBOX[13].sbox/z[9] ), .Z(n2795) );
  XOR \b/SBOX[13].sbox/U126  ( .A(\b/SBOX[13].sbox/z[1] ), .B(
        \b/SBOX[13].sbox/z[2] ), .Z(n2796) );
  XOR \b/SBOX[13].sbox/U125  ( .A(n2845), .B(n2797), .Z(shift_row_out[76]) );
  XOR \b/SBOX[13].sbox/U124  ( .A(\b/SBOX[13].sbox/z[3] ), .B(n2846), .Z(n2797) );
  XOR \b/SBOX[13].sbox/U123  ( .A(n2847), .B(n2798), .Z(shift_row_out[79]) );
  XOR \b/SBOX[13].sbox/U122  ( .A(\b/SBOX[13].sbox/z[6] ), .B(
        \b/SBOX[13].sbox/z[9] ), .Z(n2798) );
  XOR \b/SBOX[13].sbox/U121  ( .A(n2800), .B(n2799), .Z(n2848) );
  XOR \b/SBOX[13].sbox/U120  ( .A(n2802), .B(n2801), .Z(n2799) );
  XOR \b/SBOX[13].sbox/U119  ( .A(msg[109]), .B(msg[105]), .Z(n2800) );
  XOR \b/SBOX[13].sbox/U118  ( .A(\b/SBOX[13].sbox/t[36] ), .B(
        \b/SBOX[13].sbox/t[39] ), .Z(n2801) );
  XOR \b/SBOX[13].sbox/U117  ( .A(\b/SBOX[13].sbox/t[3] ), .B(
        \b/SBOX[13].sbox/t[8] ), .Z(n2802) );
  XOR \b/SBOX[13].sbox/U116  ( .A(n2804), .B(n2803), .Z(
        \b/SBOX[13].sbox/t[41] ) );
  XOR \b/SBOX[13].sbox/U115  ( .A(n2848), .B(n2805), .Z(n2803) );
  XOR \b/SBOX[13].sbox/U114  ( .A(\b/SBOX[13].sbox/t[32] ), .B(msg[111]), .Z(
        n2804) );
  XOR \b/SBOX[13].sbox/U113  ( .A(\b/SBOX[13].sbox/t[5] ), .B(
        \b/SBOX[13].sbox/t[10] ), .Z(n2805) );
  XOR \b/SBOX[13].sbox/U112  ( .A(\b/SBOX[13].sbox/t[2] ), .B(msg[110]), .Z(
        n2849) );
  XOR \b/SBOX[13].sbox/U111  ( .A(n2807), .B(n2806), .Z(
        \b/SBOX[13].sbox/t[45] ) );
  XOR \b/SBOX[13].sbox/U110  ( .A(n2849), .B(n2808), .Z(n2806) );
  XOR \b/SBOX[13].sbox/U109  ( .A(msg[108]), .B(n2848), .Z(n2807) );
  XOR \b/SBOX[13].sbox/U108  ( .A(\b/SBOX[13].sbox/t[7] ), .B(
        \b/SBOX[13].sbox/t[28] ), .Z(n2808) );
  XOR \b/SBOX[13].sbox/U107  ( .A(n2849), .B(n2809), .Z(n2854) );
  XOR \b/SBOX[13].sbox/U106  ( .A(\b/SBOX[13].sbox/t[5] ), .B(msg[108]), .Z(
        n2809) );
  XOR \b/SBOX[13].sbox/U105  ( .A(msg[111]), .B(n2810), .Z(n2850) );
  XOR \b/SBOX[13].sbox/U104  ( .A(\b/SBOX[13].sbox/t[7] ), .B(
        \b/SBOX[13].sbox/t[10] ), .Z(n2810) );
  XOR \b/SBOX[13].sbox/U103  ( .A(n2812), .B(n2811), .Z(
        \b/SBOX[13].sbox/t[42] ) );
  XOR \b/SBOX[13].sbox/U102  ( .A(n2854), .B(n2850), .Z(n2811) );
  XOR \b/SBOX[13].sbox/U101  ( .A(\b/SBOX[13].sbox/t[28] ), .B(
        \b/SBOX[13].sbox/t[32] ), .Z(n2812) );
  XOR \b/SBOX[13].sbox/U100  ( .A(msg[105]), .B(n2813), .Z(n2852) );
  XOR \b/SBOX[13].sbox/U99  ( .A(msg[107]), .B(msg[106]), .Z(n2813) );
  XOR \b/SBOX[13].sbox/U98  ( .A(msg[109]), .B(n2852), .Z(
        \b/SBOX[13].sbox/y[16] ) );
  XOR \b/SBOX[13].sbox/U97  ( .A(\b/SBOX[13].sbox/y[16] ), .B(n2814), .Z(n2853) );
  XOR \b/SBOX[13].sbox/U96  ( .A(\b/SBOX[13].sbox/t[12] ), .B(
        \b/SBOX[13].sbox/t[15] ), .Z(n2814) );
  XOR \b/SBOX[13].sbox/U95  ( .A(n2853), .B(n2815), .Z(\b/SBOX[13].sbox/t[29] ) );
  XOR \b/SBOX[13].sbox/U94  ( .A(\b/SBOX[13].sbox/t[28] ), .B(n2854), .Z(n2815) );
  XOR \b/SBOX[13].sbox/U93  ( .A(msg[104]), .B(n2816), .Z(
        \b/SBOX[13].sbox/y[1] ) );
  XOR \b/SBOX[13].sbox/U92  ( .A(msg[110]), .B(msg[109]), .Z(n2816) );
  XOR \b/SBOX[13].sbox/U91  ( .A(msg[111]), .B(\b/SBOX[13].sbox/y[1] ), .Z(
        \b/SBOX[13].sbox/y[2] ) );
  XOR \b/SBOX[13].sbox/U90  ( .A(n2818), .B(n2817), .Z(\b/SBOX[13].sbox/t[25] ) );
  XOR \b/SBOX[13].sbox/U89  ( .A(n2820), .B(n2819), .Z(n2817) );
  XOR \b/SBOX[13].sbox/U88  ( .A(msg[111]), .B(msg[109]), .Z(n2818) );
  XOR \b/SBOX[13].sbox/U87  ( .A(\b/SBOX[13].sbox/t[13] ), .B(
        \b/SBOX[13].sbox/t[15] ), .Z(n2819) );
  XOR \b/SBOX[13].sbox/U86  ( .A(\b/SBOX[13].sbox/t[3] ), .B(
        \b/SBOX[13].sbox/t[5] ), .Z(n2820) );
  XOR \b/SBOX[13].sbox/U85  ( .A(\b/SBOX[13].sbox/t[39] ), .B(
        \b/SBOX[13].sbox/t[25] ), .Z(\b/SBOX[13].sbox/t[40] ) );
  XOR \b/SBOX[13].sbox/U84  ( .A(msg[105]), .B(\b/SBOX[13].sbox/y[1] ), .Z(
        \b/SBOX[13].sbox/y[5] ) );
  XOR \b/SBOX[13].sbox/U83  ( .A(n2822), .B(n2821), .Z(\b/SBOX[13].sbox/y[15] ) );
  XOR \b/SBOX[13].sbox/U82  ( .A(msg[107]), .B(msg[105]), .Z(n2821) );
  XOR \b/SBOX[13].sbox/U81  ( .A(msg[111]), .B(msg[108]), .Z(n2822) );
  XOR \b/SBOX[13].sbox/U80  ( .A(n2824), .B(n2823), .Z(\b/SBOX[13].sbox/t[21] ) );
  XOR \b/SBOX[13].sbox/U79  ( .A(n2826), .B(n2825), .Z(n2823) );
  XOR \b/SBOX[13].sbox/U78  ( .A(\b/SBOX[13].sbox/y[15] ), .B(n2849), .Z(n2824) );
  XOR \b/SBOX[13].sbox/U77  ( .A(\b/SBOX[13].sbox/t[13] ), .B(msg[106]), .Z(
        n2825) );
  XOR \b/SBOX[13].sbox/U76  ( .A(\b/SBOX[13].sbox/t[3] ), .B(
        \b/SBOX[13].sbox/t[12] ), .Z(n2826) );
  XOR \b/SBOX[13].sbox/U75  ( .A(\b/SBOX[13].sbox/t[21] ), .B(n2827), .Z(
        \b/SBOX[13].sbox/t[43] ) );
  XOR \b/SBOX[13].sbox/U74  ( .A(\b/SBOX[13].sbox/t[28] ), .B(
        \b/SBOX[13].sbox/t[39] ), .Z(n2827) );
  XOR \b/SBOX[13].sbox/U73  ( .A(n2853), .B(n2850), .Z(\b/SBOX[13].sbox/t[24] ) );
  XOR \b/SBOX[13].sbox/U72  ( .A(\b/SBOX[13].sbox/t[32] ), .B(
        \b/SBOX[13].sbox/t[24] ), .Z(\b/SBOX[13].sbox/t[33] ) );
  XOR \b/SBOX[13].sbox/U71  ( .A(msg[108]), .B(\b/SBOX[13].sbox/y[1] ), .Z(
        \b/SBOX[13].sbox/y[4] ) );
  XOR \b/SBOX[13].sbox/U70  ( .A(n2829), .B(n2828), .Z(\b/SBOX[13].sbox/t[30] ) );
  XOR \b/SBOX[13].sbox/U69  ( .A(msg[105]), .B(n2830), .Z(n2828) );
  XOR \b/SBOX[13].sbox/U68  ( .A(\b/SBOX[13].sbox/t[13] ), .B(
        \b/SBOX[13].sbox/t[15] ), .Z(n2829) );
  XOR \b/SBOX[13].sbox/U67  ( .A(\b/SBOX[13].sbox/t[8] ), .B(
        \b/SBOX[13].sbox/t[10] ), .Z(n2830) );
  XOR \b/SBOX[13].sbox/U66  ( .A(\b/SBOX[13].sbox/t[30] ), .B(n2831), .Z(
        \b/SBOX[13].sbox/t[37] ) );
  XOR \b/SBOX[13].sbox/U65  ( .A(\b/SBOX[13].sbox/t[32] ), .B(
        \b/SBOX[13].sbox/t[36] ), .Z(n2831) );
  XOR \b/SBOX[13].sbox/U64  ( .A(msg[111]), .B(msg[106]), .Z(n2851) );
  XOR \b/SBOX[13].sbox/U63  ( .A(\b/SBOX[13].sbox/y[5] ), .B(n2851), .Z(
        \b/SBOX[13].sbox/y[3] ) );
  XOR \b/SBOX[13].sbox/U62  ( .A(n2833), .B(n2832), .Z(\b/SBOX[13].sbox/t[23] ) );
  XOR \b/SBOX[13].sbox/U61  ( .A(n2835), .B(n2834), .Z(n2832) );
  XOR \b/SBOX[13].sbox/U60  ( .A(n2851), .B(n2836), .Z(n2833) );
  XOR \b/SBOX[13].sbox/U59  ( .A(msg[109]), .B(msg[107]), .Z(n2834) );
  XOR \b/SBOX[13].sbox/U58  ( .A(\b/SBOX[13].sbox/t[12] ), .B(
        \b/SBOX[13].sbox/t[13] ), .Z(n2835) );
  XOR \b/SBOX[13].sbox/U57  ( .A(\b/SBOX[13].sbox/t[7] ), .B(
        \b/SBOX[13].sbox/t[8] ), .Z(n2836) );
  XOR \b/SBOX[13].sbox/U56  ( .A(\b/SBOX[13].sbox/t[36] ), .B(
        \b/SBOX[13].sbox/t[23] ), .Z(\b/SBOX[13].sbox/t[44] ) );
  XOR \b/SBOX[13].sbox/U55  ( .A(n2851), .B(n2837), .Z(\b/SBOX[13].sbox/y[12] ) );
  XOR \b/SBOX[13].sbox/U54  ( .A(msg[108]), .B(msg[105]), .Z(n2837) );
  XOR \b/SBOX[13].sbox/U53  ( .A(\b/SBOX[13].sbox/y[15] ), .B(n2838), .Z(
        \b/SBOX[13].sbox/y[10] ) );
  XOR \b/SBOX[13].sbox/U52  ( .A(msg[110]), .B(msg[109]), .Z(n2838) );
  XOR \b/SBOX[13].sbox/U51  ( .A(n2851), .B(n2839), .Z(\b/SBOX[13].sbox/y[17] ) );
  XOR \b/SBOX[13].sbox/U50  ( .A(msg[109]), .B(msg[108]), .Z(n2839) );
  XOR \b/SBOX[13].sbox/U49  ( .A(msg[110]), .B(n2852), .Z(
        \b/SBOX[13].sbox/y[11] ) );
  XOR \b/SBOX[13].sbox/U48  ( .A(msg[104]), .B(\b/SBOX[13].sbox/y[11] ), .Z(
        \b/SBOX[13].sbox/y[7] ) );
  XOR \b/SBOX[13].sbox/U47  ( .A(msg[104]), .B(\b/SBOX[13].sbox/y[15] ), .Z(
        \b/SBOX[13].sbox/y[6] ) );
  XOR \b/SBOX[13].sbox/U46  ( .A(\b/SBOX[13].sbox/t[26] ), .B(
        \b/SBOX[13].sbox/t[24] ), .Z(\b/SBOX[13].sbox/t[27] ) );
  XOR \b/SBOX[13].sbox/U45  ( .A(\b/SBOX[13].sbox/t[36] ), .B(
        \b/SBOX[13].sbox/t[27] ), .Z(\b/SBOX[13].sbox/t[38] ) );
  XOR \b/SBOX[13].sbox/U44  ( .A(n2853), .B(n2840), .Z(\b/SBOX[13].sbox/t[31] ) );
  XOR \b/SBOX[13].sbox/U43  ( .A(\b/SBOX[13].sbox/t[26] ), .B(n2854), .Z(n2840) );
  XOR \b/SBOX[12].sbox/U157  ( .A(\b/SBOX[12].sbox/z[12] ), .B(n2697), .Z(
        n2761) );
  XOR \b/SBOX[12].sbox/U156  ( .A(\b/SBOX[12].sbox/z[0] ), .B(
        \b/SBOX[12].sbox/z[2] ), .Z(n2697) );
  XOR \b/SBOX[12].sbox/U155  ( .A(n2699), .B(n2698), .Z(n2760) );
  XOR \b/SBOX[12].sbox/U154  ( .A(\b/SBOX[12].sbox/z[15] ), .B(
        \b/SBOX[12].sbox/z[16] ), .Z(n2698) );
  XOR \b/SBOX[12].sbox/U153  ( .A(\b/SBOX[12].sbox/z[5] ), .B(
        \b/SBOX[12].sbox/z[13] ), .Z(n2699) );
  XOR \b/SBOX[12].sbox/U152  ( .A(n2760), .B(n2700), .Z(n2774) );
  XOR \b/SBOX[12].sbox/U151  ( .A(\b/SBOX[12].sbox/z[3] ), .B(n2761), .Z(n2700) );
  XOR \b/SBOX[12].sbox/U150  ( .A(n2702), .B(n2701), .Z(n2775) );
  XOR \b/SBOX[12].sbox/U149  ( .A(n2760), .B(n2703), .Z(n2701) );
  XOR \b/SBOX[12].sbox/U148  ( .A(\b/SBOX[12].sbox/z[8] ), .B(
        \b/SBOX[12].sbox/z[12] ), .Z(n2702) );
  XOR \b/SBOX[12].sbox/U147  ( .A(\b/SBOX[12].sbox/z[4] ), .B(
        \b/SBOX[12].sbox/z[7] ), .Z(n2703) );
  XOR \b/SBOX[12].sbox/U146  ( .A(n2761), .B(n2704), .Z(n2763) );
  XOR \b/SBOX[12].sbox/U145  ( .A(\b/SBOX[12].sbox/z[8] ), .B(
        \b/SBOX[12].sbox/z[14] ), .Z(n2704) );
  XOR \b/SBOX[12].sbox/U144  ( .A(n2706), .B(n2705), .Z(n2776) );
  XOR \b/SBOX[12].sbox/U143  ( .A(\b/SBOX[12].sbox/z[17] ), .B(n2763), .Z(
        n2705) );
  XOR \b/SBOX[12].sbox/U142  ( .A(\b/SBOX[12].sbox/z[6] ), .B(
        \b/SBOX[12].sbox/z[15] ), .Z(n2706) );
  XOR \b/SBOX[12].sbox/U141  ( .A(\b/SBOX[12].sbox/z[9] ), .B(n2707), .Z(n2764) );
  XOR \b/SBOX[12].sbox/U140  ( .A(\b/SBOX[12].sbox/z[0] ), .B(
        \b/SBOX[12].sbox/z[1] ), .Z(n2707) );
  XOR \b/SBOX[12].sbox/U139  ( .A(\b/SBOX[12].sbox/z[16] ), .B(n2708), .Z(
        n2762) );
  XOR \b/SBOX[12].sbox/U138  ( .A(\b/SBOX[12].sbox/z[10] ), .B(
        \b/SBOX[12].sbox/z[15] ), .Z(n2708) );
  XOR \b/SBOX[12].sbox/U137  ( .A(n2710), .B(n2709), .Z(n2777) );
  XOR \b/SBOX[12].sbox/U136  ( .A(n2764), .B(n2762), .Z(n2709) );
  XOR \b/SBOX[12].sbox/U135  ( .A(\b/SBOX[12].sbox/z[6] ), .B(
        \b/SBOX[12].sbox/z[7] ), .Z(n2710) );
  XOR \b/SBOX[12].sbox/U134  ( .A(\b/SBOX[12].sbox/z[4] ), .B(n2762), .Z(n2765) );
  XOR \b/SBOX[12].sbox/U133  ( .A(n2765), .B(n2711), .Z(n2766) );
  XOR \b/SBOX[12].sbox/U132  ( .A(\b/SBOX[12].sbox/z[3] ), .B(
        \b/SBOX[12].sbox/z[7] ), .Z(n2711) );
  XOR \b/SBOX[12].sbox/U131  ( .A(n2763), .B(n2712), .Z(shift_row_out[98]) );
  XOR \b/SBOX[12].sbox/U130  ( .A(\b/SBOX[12].sbox/z[11] ), .B(n2766), .Z(
        n2712) );
  XOR \b/SBOX[12].sbox/U129  ( .A(n2714), .B(n2713), .Z(shift_row_out[99]) );
  XOR \b/SBOX[12].sbox/U128  ( .A(n2765), .B(n2715), .Z(n2713) );
  XOR \b/SBOX[12].sbox/U127  ( .A(\b/SBOX[12].sbox/z[5] ), .B(
        \b/SBOX[12].sbox/z[9] ), .Z(n2714) );
  XOR \b/SBOX[12].sbox/U126  ( .A(\b/SBOX[12].sbox/z[1] ), .B(
        \b/SBOX[12].sbox/z[2] ), .Z(n2715) );
  XOR \b/SBOX[12].sbox/U125  ( .A(n2764), .B(n2716), .Z(shift_row_out[100]) );
  XOR \b/SBOX[12].sbox/U124  ( .A(\b/SBOX[12].sbox/z[3] ), .B(n2765), .Z(n2716) );
  XOR \b/SBOX[12].sbox/U123  ( .A(n2766), .B(n2717), .Z(shift_row_out[103]) );
  XOR \b/SBOX[12].sbox/U122  ( .A(\b/SBOX[12].sbox/z[6] ), .B(
        \b/SBOX[12].sbox/z[9] ), .Z(n2717) );
  XOR \b/SBOX[12].sbox/U121  ( .A(n2719), .B(n2718), .Z(n2767) );
  XOR \b/SBOX[12].sbox/U120  ( .A(n2721), .B(n2720), .Z(n2718) );
  XOR \b/SBOX[12].sbox/U119  ( .A(msg[101]), .B(msg[97]), .Z(n2719) );
  XOR \b/SBOX[12].sbox/U118  ( .A(\b/SBOX[12].sbox/t[36] ), .B(
        \b/SBOX[12].sbox/t[39] ), .Z(n2720) );
  XOR \b/SBOX[12].sbox/U117  ( .A(\b/SBOX[12].sbox/t[3] ), .B(
        \b/SBOX[12].sbox/t[8] ), .Z(n2721) );
  XOR \b/SBOX[12].sbox/U116  ( .A(n2723), .B(n2722), .Z(
        \b/SBOX[12].sbox/t[41] ) );
  XOR \b/SBOX[12].sbox/U115  ( .A(n2767), .B(n2724), .Z(n2722) );
  XOR \b/SBOX[12].sbox/U114  ( .A(\b/SBOX[12].sbox/t[32] ), .B(msg[103]), .Z(
        n2723) );
  XOR \b/SBOX[12].sbox/U113  ( .A(\b/SBOX[12].sbox/t[5] ), .B(
        \b/SBOX[12].sbox/t[10] ), .Z(n2724) );
  XOR \b/SBOX[12].sbox/U112  ( .A(\b/SBOX[12].sbox/t[2] ), .B(msg[102]), .Z(
        n2768) );
  XOR \b/SBOX[12].sbox/U111  ( .A(n2726), .B(n2725), .Z(
        \b/SBOX[12].sbox/t[45] ) );
  XOR \b/SBOX[12].sbox/U110  ( .A(n2768), .B(n2727), .Z(n2725) );
  XOR \b/SBOX[12].sbox/U109  ( .A(msg[100]), .B(n2767), .Z(n2726) );
  XOR \b/SBOX[12].sbox/U108  ( .A(\b/SBOX[12].sbox/t[7] ), .B(
        \b/SBOX[12].sbox/t[28] ), .Z(n2727) );
  XOR \b/SBOX[12].sbox/U107  ( .A(n2768), .B(n2728), .Z(n2773) );
  XOR \b/SBOX[12].sbox/U106  ( .A(\b/SBOX[12].sbox/t[5] ), .B(msg[100]), .Z(
        n2728) );
  XOR \b/SBOX[12].sbox/U105  ( .A(msg[103]), .B(n2729), .Z(n2769) );
  XOR \b/SBOX[12].sbox/U104  ( .A(\b/SBOX[12].sbox/t[7] ), .B(
        \b/SBOX[12].sbox/t[10] ), .Z(n2729) );
  XOR \b/SBOX[12].sbox/U103  ( .A(n2731), .B(n2730), .Z(
        \b/SBOX[12].sbox/t[42] ) );
  XOR \b/SBOX[12].sbox/U102  ( .A(n2773), .B(n2769), .Z(n2730) );
  XOR \b/SBOX[12].sbox/U101  ( .A(\b/SBOX[12].sbox/t[28] ), .B(
        \b/SBOX[12].sbox/t[32] ), .Z(n2731) );
  XOR \b/SBOX[12].sbox/U100  ( .A(msg[97]), .B(n2732), .Z(n2771) );
  XOR \b/SBOX[12].sbox/U99  ( .A(msg[99]), .B(msg[98]), .Z(n2732) );
  XOR \b/SBOX[12].sbox/U98  ( .A(msg[101]), .B(n2771), .Z(
        \b/SBOX[12].sbox/y[16] ) );
  XOR \b/SBOX[12].sbox/U97  ( .A(\b/SBOX[12].sbox/y[16] ), .B(n2733), .Z(n2772) );
  XOR \b/SBOX[12].sbox/U96  ( .A(\b/SBOX[12].sbox/t[12] ), .B(
        \b/SBOX[12].sbox/t[15] ), .Z(n2733) );
  XOR \b/SBOX[12].sbox/U95  ( .A(n2772), .B(n2734), .Z(\b/SBOX[12].sbox/t[29] ) );
  XOR \b/SBOX[12].sbox/U94  ( .A(\b/SBOX[12].sbox/t[28] ), .B(n2773), .Z(n2734) );
  XOR \b/SBOX[12].sbox/U93  ( .A(msg[96]), .B(n2735), .Z(
        \b/SBOX[12].sbox/y[1] ) );
  XOR \b/SBOX[12].sbox/U92  ( .A(msg[102]), .B(msg[101]), .Z(n2735) );
  XOR \b/SBOX[12].sbox/U91  ( .A(msg[103]), .B(\b/SBOX[12].sbox/y[1] ), .Z(
        \b/SBOX[12].sbox/y[2] ) );
  XOR \b/SBOX[12].sbox/U90  ( .A(n2737), .B(n2736), .Z(\b/SBOX[12].sbox/t[25] ) );
  XOR \b/SBOX[12].sbox/U89  ( .A(n2739), .B(n2738), .Z(n2736) );
  XOR \b/SBOX[12].sbox/U88  ( .A(msg[103]), .B(msg[101]), .Z(n2737) );
  XOR \b/SBOX[12].sbox/U87  ( .A(\b/SBOX[12].sbox/t[13] ), .B(
        \b/SBOX[12].sbox/t[15] ), .Z(n2738) );
  XOR \b/SBOX[12].sbox/U86  ( .A(\b/SBOX[12].sbox/t[3] ), .B(
        \b/SBOX[12].sbox/t[5] ), .Z(n2739) );
  XOR \b/SBOX[12].sbox/U85  ( .A(\b/SBOX[12].sbox/t[39] ), .B(
        \b/SBOX[12].sbox/t[25] ), .Z(\b/SBOX[12].sbox/t[40] ) );
  XOR \b/SBOX[12].sbox/U84  ( .A(msg[97]), .B(\b/SBOX[12].sbox/y[1] ), .Z(
        \b/SBOX[12].sbox/y[5] ) );
  XOR \b/SBOX[12].sbox/U83  ( .A(n2741), .B(n2740), .Z(\b/SBOX[12].sbox/y[15] ) );
  XOR \b/SBOX[12].sbox/U82  ( .A(msg[99]), .B(msg[97]), .Z(n2740) );
  XOR \b/SBOX[12].sbox/U81  ( .A(msg[103]), .B(msg[100]), .Z(n2741) );
  XOR \b/SBOX[12].sbox/U80  ( .A(n2743), .B(n2742), .Z(\b/SBOX[12].sbox/t[21] ) );
  XOR \b/SBOX[12].sbox/U79  ( .A(n2745), .B(n2744), .Z(n2742) );
  XOR \b/SBOX[12].sbox/U78  ( .A(\b/SBOX[12].sbox/y[15] ), .B(n2768), .Z(n2743) );
  XOR \b/SBOX[12].sbox/U77  ( .A(\b/SBOX[12].sbox/t[13] ), .B(msg[98]), .Z(
        n2744) );
  XOR \b/SBOX[12].sbox/U76  ( .A(\b/SBOX[12].sbox/t[3] ), .B(
        \b/SBOX[12].sbox/t[12] ), .Z(n2745) );
  XOR \b/SBOX[12].sbox/U75  ( .A(\b/SBOX[12].sbox/t[21] ), .B(n2746), .Z(
        \b/SBOX[12].sbox/t[43] ) );
  XOR \b/SBOX[12].sbox/U74  ( .A(\b/SBOX[12].sbox/t[28] ), .B(
        \b/SBOX[12].sbox/t[39] ), .Z(n2746) );
  XOR \b/SBOX[12].sbox/U73  ( .A(n2772), .B(n2769), .Z(\b/SBOX[12].sbox/t[24] ) );
  XOR \b/SBOX[12].sbox/U72  ( .A(\b/SBOX[12].sbox/t[32] ), .B(
        \b/SBOX[12].sbox/t[24] ), .Z(\b/SBOX[12].sbox/t[33] ) );
  XOR \b/SBOX[12].sbox/U71  ( .A(msg[100]), .B(\b/SBOX[12].sbox/y[1] ), .Z(
        \b/SBOX[12].sbox/y[4] ) );
  XOR \b/SBOX[12].sbox/U70  ( .A(n2748), .B(n2747), .Z(\b/SBOX[12].sbox/t[30] ) );
  XOR \b/SBOX[12].sbox/U69  ( .A(msg[97]), .B(n2749), .Z(n2747) );
  XOR \b/SBOX[12].sbox/U68  ( .A(\b/SBOX[12].sbox/t[13] ), .B(
        \b/SBOX[12].sbox/t[15] ), .Z(n2748) );
  XOR \b/SBOX[12].sbox/U67  ( .A(\b/SBOX[12].sbox/t[8] ), .B(
        \b/SBOX[12].sbox/t[10] ), .Z(n2749) );
  XOR \b/SBOX[12].sbox/U66  ( .A(\b/SBOX[12].sbox/t[30] ), .B(n2750), .Z(
        \b/SBOX[12].sbox/t[37] ) );
  XOR \b/SBOX[12].sbox/U65  ( .A(\b/SBOX[12].sbox/t[32] ), .B(
        \b/SBOX[12].sbox/t[36] ), .Z(n2750) );
  XOR \b/SBOX[12].sbox/U64  ( .A(msg[103]), .B(msg[98]), .Z(n2770) );
  XOR \b/SBOX[12].sbox/U63  ( .A(\b/SBOX[12].sbox/y[5] ), .B(n2770), .Z(
        \b/SBOX[12].sbox/y[3] ) );
  XOR \b/SBOX[12].sbox/U62  ( .A(n2752), .B(n2751), .Z(\b/SBOX[12].sbox/t[23] ) );
  XOR \b/SBOX[12].sbox/U61  ( .A(n2754), .B(n2753), .Z(n2751) );
  XOR \b/SBOX[12].sbox/U60  ( .A(n2770), .B(n2755), .Z(n2752) );
  XOR \b/SBOX[12].sbox/U59  ( .A(msg[101]), .B(msg[99]), .Z(n2753) );
  XOR \b/SBOX[12].sbox/U58  ( .A(\b/SBOX[12].sbox/t[12] ), .B(
        \b/SBOX[12].sbox/t[13] ), .Z(n2754) );
  XOR \b/SBOX[12].sbox/U57  ( .A(\b/SBOX[12].sbox/t[7] ), .B(
        \b/SBOX[12].sbox/t[8] ), .Z(n2755) );
  XOR \b/SBOX[12].sbox/U56  ( .A(\b/SBOX[12].sbox/t[36] ), .B(
        \b/SBOX[12].sbox/t[23] ), .Z(\b/SBOX[12].sbox/t[44] ) );
  XOR \b/SBOX[12].sbox/U55  ( .A(n2770), .B(n2756), .Z(\b/SBOX[12].sbox/y[12] ) );
  XOR \b/SBOX[12].sbox/U54  ( .A(msg[100]), .B(msg[97]), .Z(n2756) );
  XOR \b/SBOX[12].sbox/U53  ( .A(\b/SBOX[12].sbox/y[15] ), .B(n2757), .Z(
        \b/SBOX[12].sbox/y[10] ) );
  XOR \b/SBOX[12].sbox/U52  ( .A(msg[102]), .B(msg[101]), .Z(n2757) );
  XOR \b/SBOX[12].sbox/U51  ( .A(n2770), .B(n2758), .Z(\b/SBOX[12].sbox/y[17] ) );
  XOR \b/SBOX[12].sbox/U50  ( .A(msg[101]), .B(msg[100]), .Z(n2758) );
  XOR \b/SBOX[12].sbox/U49  ( .A(msg[102]), .B(n2771), .Z(
        \b/SBOX[12].sbox/y[11] ) );
  XOR \b/SBOX[12].sbox/U48  ( .A(msg[96]), .B(\b/SBOX[12].sbox/y[11] ), .Z(
        \b/SBOX[12].sbox/y[7] ) );
  XOR \b/SBOX[12].sbox/U47  ( .A(msg[96]), .B(\b/SBOX[12].sbox/y[15] ), .Z(
        \b/SBOX[12].sbox/y[6] ) );
  XOR \b/SBOX[12].sbox/U46  ( .A(\b/SBOX[12].sbox/t[26] ), .B(
        \b/SBOX[12].sbox/t[24] ), .Z(\b/SBOX[12].sbox/t[27] ) );
  XOR \b/SBOX[12].sbox/U45  ( .A(\b/SBOX[12].sbox/t[36] ), .B(
        \b/SBOX[12].sbox/t[27] ), .Z(\b/SBOX[12].sbox/t[38] ) );
  XOR \b/SBOX[12].sbox/U44  ( .A(n2772), .B(n2759), .Z(\b/SBOX[12].sbox/t[31] ) );
  XOR \b/SBOX[12].sbox/U43  ( .A(\b/SBOX[12].sbox/t[26] ), .B(n2773), .Z(n2759) );
  XOR \b/SBOX[11].sbox/U157  ( .A(\b/SBOX[11].sbox/z[12] ), .B(n2616), .Z(
        n2680) );
  XOR \b/SBOX[11].sbox/U156  ( .A(\b/SBOX[11].sbox/z[0] ), .B(
        \b/SBOX[11].sbox/z[2] ), .Z(n2616) );
  XOR \b/SBOX[11].sbox/U155  ( .A(n2618), .B(n2617), .Z(n2679) );
  XOR \b/SBOX[11].sbox/U154  ( .A(\b/SBOX[11].sbox/z[15] ), .B(
        \b/SBOX[11].sbox/z[16] ), .Z(n2617) );
  XOR \b/SBOX[11].sbox/U153  ( .A(\b/SBOX[11].sbox/z[5] ), .B(
        \b/SBOX[11].sbox/z[13] ), .Z(n2618) );
  XOR \b/SBOX[11].sbox/U152  ( .A(n2679), .B(n2619), .Z(n2693) );
  XOR \b/SBOX[11].sbox/U151  ( .A(\b/SBOX[11].sbox/z[3] ), .B(n2680), .Z(n2619) );
  XOR \b/SBOX[11].sbox/U150  ( .A(n2621), .B(n2620), .Z(n2694) );
  XOR \b/SBOX[11].sbox/U149  ( .A(n2679), .B(n2622), .Z(n2620) );
  XOR \b/SBOX[11].sbox/U148  ( .A(\b/SBOX[11].sbox/z[8] ), .B(
        \b/SBOX[11].sbox/z[12] ), .Z(n2621) );
  XOR \b/SBOX[11].sbox/U147  ( .A(\b/SBOX[11].sbox/z[4] ), .B(
        \b/SBOX[11].sbox/z[7] ), .Z(n2622) );
  XOR \b/SBOX[11].sbox/U146  ( .A(n2680), .B(n2623), .Z(n2682) );
  XOR \b/SBOX[11].sbox/U145  ( .A(\b/SBOX[11].sbox/z[8] ), .B(
        \b/SBOX[11].sbox/z[14] ), .Z(n2623) );
  XOR \b/SBOX[11].sbox/U144  ( .A(n2625), .B(n2624), .Z(n2695) );
  XOR \b/SBOX[11].sbox/U143  ( .A(\b/SBOX[11].sbox/z[17] ), .B(n2682), .Z(
        n2624) );
  XOR \b/SBOX[11].sbox/U142  ( .A(\b/SBOX[11].sbox/z[6] ), .B(
        \b/SBOX[11].sbox/z[15] ), .Z(n2625) );
  XOR \b/SBOX[11].sbox/U141  ( .A(\b/SBOX[11].sbox/z[9] ), .B(n2626), .Z(n2683) );
  XOR \b/SBOX[11].sbox/U140  ( .A(\b/SBOX[11].sbox/z[0] ), .B(
        \b/SBOX[11].sbox/z[1] ), .Z(n2626) );
  XOR \b/SBOX[11].sbox/U139  ( .A(\b/SBOX[11].sbox/z[16] ), .B(n2627), .Z(
        n2681) );
  XOR \b/SBOX[11].sbox/U138  ( .A(\b/SBOX[11].sbox/z[10] ), .B(
        \b/SBOX[11].sbox/z[15] ), .Z(n2627) );
  XOR \b/SBOX[11].sbox/U137  ( .A(n2629), .B(n2628), .Z(n2696) );
  XOR \b/SBOX[11].sbox/U136  ( .A(n2683), .B(n2681), .Z(n2628) );
  XOR \b/SBOX[11].sbox/U135  ( .A(\b/SBOX[11].sbox/z[6] ), .B(
        \b/SBOX[11].sbox/z[7] ), .Z(n2629) );
  XOR \b/SBOX[11].sbox/U134  ( .A(\b/SBOX[11].sbox/z[4] ), .B(n2681), .Z(n2684) );
  XOR \b/SBOX[11].sbox/U133  ( .A(n2684), .B(n2630), .Z(n2685) );
  XOR \b/SBOX[11].sbox/U132  ( .A(\b/SBOX[11].sbox/z[3] ), .B(
        \b/SBOX[11].sbox/z[7] ), .Z(n2630) );
  XOR \b/SBOX[11].sbox/U131  ( .A(n2682), .B(n2631), .Z(shift_row_out[122]) );
  XOR \b/SBOX[11].sbox/U130  ( .A(\b/SBOX[11].sbox/z[11] ), .B(n2685), .Z(
        n2631) );
  XOR \b/SBOX[11].sbox/U129  ( .A(n2633), .B(n2632), .Z(shift_row_out[123]) );
  XOR \b/SBOX[11].sbox/U128  ( .A(n2684), .B(n2634), .Z(n2632) );
  XOR \b/SBOX[11].sbox/U127  ( .A(\b/SBOX[11].sbox/z[5] ), .B(
        \b/SBOX[11].sbox/z[9] ), .Z(n2633) );
  XOR \b/SBOX[11].sbox/U126  ( .A(\b/SBOX[11].sbox/z[1] ), .B(
        \b/SBOX[11].sbox/z[2] ), .Z(n2634) );
  XOR \b/SBOX[11].sbox/U125  ( .A(n2683), .B(n2635), .Z(shift_row_out[124]) );
  XOR \b/SBOX[11].sbox/U124  ( .A(\b/SBOX[11].sbox/z[3] ), .B(n2684), .Z(n2635) );
  XOR \b/SBOX[11].sbox/U123  ( .A(n2685), .B(n2636), .Z(shift_row_out[127]) );
  XOR \b/SBOX[11].sbox/U122  ( .A(\b/SBOX[11].sbox/z[6] ), .B(
        \b/SBOX[11].sbox/z[9] ), .Z(n2636) );
  XOR \b/SBOX[11].sbox/U121  ( .A(n2638), .B(n2637), .Z(n2686) );
  XOR \b/SBOX[11].sbox/U120  ( .A(n2640), .B(n2639), .Z(n2637) );
  XOR \b/SBOX[11].sbox/U119  ( .A(msg[93]), .B(msg[89]), .Z(n2638) );
  XOR \b/SBOX[11].sbox/U118  ( .A(\b/SBOX[11].sbox/t[36] ), .B(
        \b/SBOX[11].sbox/t[39] ), .Z(n2639) );
  XOR \b/SBOX[11].sbox/U117  ( .A(\b/SBOX[11].sbox/t[3] ), .B(
        \b/SBOX[11].sbox/t[8] ), .Z(n2640) );
  XOR \b/SBOX[11].sbox/U116  ( .A(n2642), .B(n2641), .Z(
        \b/SBOX[11].sbox/t[41] ) );
  XOR \b/SBOX[11].sbox/U115  ( .A(n2686), .B(n2643), .Z(n2641) );
  XOR \b/SBOX[11].sbox/U114  ( .A(\b/SBOX[11].sbox/t[32] ), .B(msg[95]), .Z(
        n2642) );
  XOR \b/SBOX[11].sbox/U113  ( .A(\b/SBOX[11].sbox/t[5] ), .B(
        \b/SBOX[11].sbox/t[10] ), .Z(n2643) );
  XOR \b/SBOX[11].sbox/U112  ( .A(\b/SBOX[11].sbox/t[2] ), .B(msg[94]), .Z(
        n2687) );
  XOR \b/SBOX[11].sbox/U111  ( .A(n2645), .B(n2644), .Z(
        \b/SBOX[11].sbox/t[45] ) );
  XOR \b/SBOX[11].sbox/U110  ( .A(n2687), .B(n2646), .Z(n2644) );
  XOR \b/SBOX[11].sbox/U109  ( .A(msg[92]), .B(n2686), .Z(n2645) );
  XOR \b/SBOX[11].sbox/U108  ( .A(\b/SBOX[11].sbox/t[7] ), .B(
        \b/SBOX[11].sbox/t[28] ), .Z(n2646) );
  XOR \b/SBOX[11].sbox/U107  ( .A(n2687), .B(n2647), .Z(n2692) );
  XOR \b/SBOX[11].sbox/U106  ( .A(\b/SBOX[11].sbox/t[5] ), .B(msg[92]), .Z(
        n2647) );
  XOR \b/SBOX[11].sbox/U105  ( .A(msg[95]), .B(n2648), .Z(n2688) );
  XOR \b/SBOX[11].sbox/U104  ( .A(\b/SBOX[11].sbox/t[7] ), .B(
        \b/SBOX[11].sbox/t[10] ), .Z(n2648) );
  XOR \b/SBOX[11].sbox/U103  ( .A(n2650), .B(n2649), .Z(
        \b/SBOX[11].sbox/t[42] ) );
  XOR \b/SBOX[11].sbox/U102  ( .A(n2692), .B(n2688), .Z(n2649) );
  XOR \b/SBOX[11].sbox/U101  ( .A(\b/SBOX[11].sbox/t[28] ), .B(
        \b/SBOX[11].sbox/t[32] ), .Z(n2650) );
  XOR \b/SBOX[11].sbox/U100  ( .A(msg[89]), .B(n2651), .Z(n2690) );
  XOR \b/SBOX[11].sbox/U99  ( .A(msg[91]), .B(msg[90]), .Z(n2651) );
  XOR \b/SBOX[11].sbox/U98  ( .A(msg[93]), .B(n2690), .Z(
        \b/SBOX[11].sbox/y[16] ) );
  XOR \b/SBOX[11].sbox/U97  ( .A(\b/SBOX[11].sbox/y[16] ), .B(n2652), .Z(n2691) );
  XOR \b/SBOX[11].sbox/U96  ( .A(\b/SBOX[11].sbox/t[12] ), .B(
        \b/SBOX[11].sbox/t[15] ), .Z(n2652) );
  XOR \b/SBOX[11].sbox/U95  ( .A(n2691), .B(n2653), .Z(\b/SBOX[11].sbox/t[29] ) );
  XOR \b/SBOX[11].sbox/U94  ( .A(\b/SBOX[11].sbox/t[28] ), .B(n2692), .Z(n2653) );
  XOR \b/SBOX[11].sbox/U93  ( .A(msg[88]), .B(n2654), .Z(
        \b/SBOX[11].sbox/y[1] ) );
  XOR \b/SBOX[11].sbox/U92  ( .A(msg[94]), .B(msg[93]), .Z(n2654) );
  XOR \b/SBOX[11].sbox/U91  ( .A(msg[95]), .B(\b/SBOX[11].sbox/y[1] ), .Z(
        \b/SBOX[11].sbox/y[2] ) );
  XOR \b/SBOX[11].sbox/U90  ( .A(n2656), .B(n2655), .Z(\b/SBOX[11].sbox/t[25] ) );
  XOR \b/SBOX[11].sbox/U89  ( .A(n2658), .B(n2657), .Z(n2655) );
  XOR \b/SBOX[11].sbox/U88  ( .A(msg[95]), .B(msg[93]), .Z(n2656) );
  XOR \b/SBOX[11].sbox/U87  ( .A(\b/SBOX[11].sbox/t[13] ), .B(
        \b/SBOX[11].sbox/t[15] ), .Z(n2657) );
  XOR \b/SBOX[11].sbox/U86  ( .A(\b/SBOX[11].sbox/t[3] ), .B(
        \b/SBOX[11].sbox/t[5] ), .Z(n2658) );
  XOR \b/SBOX[11].sbox/U85  ( .A(\b/SBOX[11].sbox/t[39] ), .B(
        \b/SBOX[11].sbox/t[25] ), .Z(\b/SBOX[11].sbox/t[40] ) );
  XOR \b/SBOX[11].sbox/U84  ( .A(msg[89]), .B(\b/SBOX[11].sbox/y[1] ), .Z(
        \b/SBOX[11].sbox/y[5] ) );
  XOR \b/SBOX[11].sbox/U83  ( .A(n2660), .B(n2659), .Z(\b/SBOX[11].sbox/y[15] ) );
  XOR \b/SBOX[11].sbox/U82  ( .A(msg[91]), .B(msg[89]), .Z(n2659) );
  XOR \b/SBOX[11].sbox/U81  ( .A(msg[95]), .B(msg[92]), .Z(n2660) );
  XOR \b/SBOX[11].sbox/U80  ( .A(n2662), .B(n2661), .Z(\b/SBOX[11].sbox/t[21] ) );
  XOR \b/SBOX[11].sbox/U79  ( .A(n2664), .B(n2663), .Z(n2661) );
  XOR \b/SBOX[11].sbox/U78  ( .A(\b/SBOX[11].sbox/y[15] ), .B(n2687), .Z(n2662) );
  XOR \b/SBOX[11].sbox/U77  ( .A(\b/SBOX[11].sbox/t[13] ), .B(msg[90]), .Z(
        n2663) );
  XOR \b/SBOX[11].sbox/U76  ( .A(\b/SBOX[11].sbox/t[3] ), .B(
        \b/SBOX[11].sbox/t[12] ), .Z(n2664) );
  XOR \b/SBOX[11].sbox/U75  ( .A(\b/SBOX[11].sbox/t[21] ), .B(n2665), .Z(
        \b/SBOX[11].sbox/t[43] ) );
  XOR \b/SBOX[11].sbox/U74  ( .A(\b/SBOX[11].sbox/t[28] ), .B(
        \b/SBOX[11].sbox/t[39] ), .Z(n2665) );
  XOR \b/SBOX[11].sbox/U73  ( .A(n2691), .B(n2688), .Z(\b/SBOX[11].sbox/t[24] ) );
  XOR \b/SBOX[11].sbox/U72  ( .A(\b/SBOX[11].sbox/t[32] ), .B(
        \b/SBOX[11].sbox/t[24] ), .Z(\b/SBOX[11].sbox/t[33] ) );
  XOR \b/SBOX[11].sbox/U71  ( .A(msg[92]), .B(\b/SBOX[11].sbox/y[1] ), .Z(
        \b/SBOX[11].sbox/y[4] ) );
  XOR \b/SBOX[11].sbox/U70  ( .A(n2667), .B(n2666), .Z(\b/SBOX[11].sbox/t[30] ) );
  XOR \b/SBOX[11].sbox/U69  ( .A(msg[89]), .B(n2668), .Z(n2666) );
  XOR \b/SBOX[11].sbox/U68  ( .A(\b/SBOX[11].sbox/t[13] ), .B(
        \b/SBOX[11].sbox/t[15] ), .Z(n2667) );
  XOR \b/SBOX[11].sbox/U67  ( .A(\b/SBOX[11].sbox/t[8] ), .B(
        \b/SBOX[11].sbox/t[10] ), .Z(n2668) );
  XOR \b/SBOX[11].sbox/U66  ( .A(\b/SBOX[11].sbox/t[30] ), .B(n2669), .Z(
        \b/SBOX[11].sbox/t[37] ) );
  XOR \b/SBOX[11].sbox/U65  ( .A(\b/SBOX[11].sbox/t[32] ), .B(
        \b/SBOX[11].sbox/t[36] ), .Z(n2669) );
  XOR \b/SBOX[11].sbox/U64  ( .A(msg[95]), .B(msg[90]), .Z(n2689) );
  XOR \b/SBOX[11].sbox/U63  ( .A(\b/SBOX[11].sbox/y[5] ), .B(n2689), .Z(
        \b/SBOX[11].sbox/y[3] ) );
  XOR \b/SBOX[11].sbox/U62  ( .A(n2671), .B(n2670), .Z(\b/SBOX[11].sbox/t[23] ) );
  XOR \b/SBOX[11].sbox/U61  ( .A(n2673), .B(n2672), .Z(n2670) );
  XOR \b/SBOX[11].sbox/U60  ( .A(n2689), .B(n2674), .Z(n2671) );
  XOR \b/SBOX[11].sbox/U59  ( .A(msg[93]), .B(msg[91]), .Z(n2672) );
  XOR \b/SBOX[11].sbox/U58  ( .A(\b/SBOX[11].sbox/t[12] ), .B(
        \b/SBOX[11].sbox/t[13] ), .Z(n2673) );
  XOR \b/SBOX[11].sbox/U57  ( .A(\b/SBOX[11].sbox/t[7] ), .B(
        \b/SBOX[11].sbox/t[8] ), .Z(n2674) );
  XOR \b/SBOX[11].sbox/U56  ( .A(\b/SBOX[11].sbox/t[36] ), .B(
        \b/SBOX[11].sbox/t[23] ), .Z(\b/SBOX[11].sbox/t[44] ) );
  XOR \b/SBOX[11].sbox/U55  ( .A(n2689), .B(n2675), .Z(\b/SBOX[11].sbox/y[12] ) );
  XOR \b/SBOX[11].sbox/U54  ( .A(msg[92]), .B(msg[89]), .Z(n2675) );
  XOR \b/SBOX[11].sbox/U53  ( .A(\b/SBOX[11].sbox/y[15] ), .B(n2676), .Z(
        \b/SBOX[11].sbox/y[10] ) );
  XOR \b/SBOX[11].sbox/U52  ( .A(msg[94]), .B(msg[93]), .Z(n2676) );
  XOR \b/SBOX[11].sbox/U51  ( .A(n2689), .B(n2677), .Z(\b/SBOX[11].sbox/y[17] ) );
  XOR \b/SBOX[11].sbox/U50  ( .A(msg[93]), .B(msg[92]), .Z(n2677) );
  XOR \b/SBOX[11].sbox/U49  ( .A(msg[94]), .B(n2690), .Z(
        \b/SBOX[11].sbox/y[11] ) );
  XOR \b/SBOX[11].sbox/U48  ( .A(msg[88]), .B(\b/SBOX[11].sbox/y[11] ), .Z(
        \b/SBOX[11].sbox/y[7] ) );
  XOR \b/SBOX[11].sbox/U47  ( .A(msg[88]), .B(\b/SBOX[11].sbox/y[15] ), .Z(
        \b/SBOX[11].sbox/y[6] ) );
  XOR \b/SBOX[11].sbox/U46  ( .A(\b/SBOX[11].sbox/t[26] ), .B(
        \b/SBOX[11].sbox/t[24] ), .Z(\b/SBOX[11].sbox/t[27] ) );
  XOR \b/SBOX[11].sbox/U45  ( .A(\b/SBOX[11].sbox/t[36] ), .B(
        \b/SBOX[11].sbox/t[27] ), .Z(\b/SBOX[11].sbox/t[38] ) );
  XOR \b/SBOX[11].sbox/U44  ( .A(n2691), .B(n2678), .Z(\b/SBOX[11].sbox/t[31] ) );
  XOR \b/SBOX[11].sbox/U43  ( .A(\b/SBOX[11].sbox/t[26] ), .B(n2692), .Z(n2678) );
  XOR \b/SBOX[10].sbox/U157  ( .A(\b/SBOX[10].sbox/z[12] ), .B(n2535), .Z(
        n2599) );
  XOR \b/SBOX[10].sbox/U156  ( .A(\b/SBOX[10].sbox/z[0] ), .B(
        \b/SBOX[10].sbox/z[2] ), .Z(n2535) );
  XOR \b/SBOX[10].sbox/U155  ( .A(n2537), .B(n2536), .Z(n2598) );
  XOR \b/SBOX[10].sbox/U154  ( .A(\b/SBOX[10].sbox/z[15] ), .B(
        \b/SBOX[10].sbox/z[16] ), .Z(n2536) );
  XOR \b/SBOX[10].sbox/U153  ( .A(\b/SBOX[10].sbox/z[5] ), .B(
        \b/SBOX[10].sbox/z[13] ), .Z(n2537) );
  XOR \b/SBOX[10].sbox/U152  ( .A(n2598), .B(n2538), .Z(n2612) );
  XOR \b/SBOX[10].sbox/U151  ( .A(\b/SBOX[10].sbox/z[3] ), .B(n2599), .Z(n2538) );
  XOR \b/SBOX[10].sbox/U150  ( .A(n2540), .B(n2539), .Z(n2613) );
  XOR \b/SBOX[10].sbox/U149  ( .A(n2598), .B(n2541), .Z(n2539) );
  XOR \b/SBOX[10].sbox/U148  ( .A(\b/SBOX[10].sbox/z[8] ), .B(
        \b/SBOX[10].sbox/z[12] ), .Z(n2540) );
  XOR \b/SBOX[10].sbox/U147  ( .A(\b/SBOX[10].sbox/z[4] ), .B(
        \b/SBOX[10].sbox/z[7] ), .Z(n2541) );
  XOR \b/SBOX[10].sbox/U146  ( .A(n2599), .B(n2542), .Z(n2601) );
  XOR \b/SBOX[10].sbox/U145  ( .A(\b/SBOX[10].sbox/z[8] ), .B(
        \b/SBOX[10].sbox/z[14] ), .Z(n2542) );
  XOR \b/SBOX[10].sbox/U144  ( .A(n2544), .B(n2543), .Z(n2614) );
  XOR \b/SBOX[10].sbox/U143  ( .A(\b/SBOX[10].sbox/z[17] ), .B(n2601), .Z(
        n2543) );
  XOR \b/SBOX[10].sbox/U142  ( .A(\b/SBOX[10].sbox/z[6] ), .B(
        \b/SBOX[10].sbox/z[15] ), .Z(n2544) );
  XOR \b/SBOX[10].sbox/U141  ( .A(\b/SBOX[10].sbox/z[9] ), .B(n2545), .Z(n2602) );
  XOR \b/SBOX[10].sbox/U140  ( .A(\b/SBOX[10].sbox/z[0] ), .B(
        \b/SBOX[10].sbox/z[1] ), .Z(n2545) );
  XOR \b/SBOX[10].sbox/U139  ( .A(\b/SBOX[10].sbox/z[16] ), .B(n2546), .Z(
        n2600) );
  XOR \b/SBOX[10].sbox/U138  ( .A(\b/SBOX[10].sbox/z[10] ), .B(
        \b/SBOX[10].sbox/z[15] ), .Z(n2546) );
  XOR \b/SBOX[10].sbox/U137  ( .A(n2548), .B(n2547), .Z(n2615) );
  XOR \b/SBOX[10].sbox/U136  ( .A(n2602), .B(n2600), .Z(n2547) );
  XOR \b/SBOX[10].sbox/U135  ( .A(\b/SBOX[10].sbox/z[6] ), .B(
        \b/SBOX[10].sbox/z[7] ), .Z(n2548) );
  XOR \b/SBOX[10].sbox/U134  ( .A(\b/SBOX[10].sbox/z[4] ), .B(n2600), .Z(n2603) );
  XOR \b/SBOX[10].sbox/U133  ( .A(n2603), .B(n2549), .Z(n2604) );
  XOR \b/SBOX[10].sbox/U132  ( .A(\b/SBOX[10].sbox/z[3] ), .B(
        \b/SBOX[10].sbox/z[7] ), .Z(n2549) );
  XOR \b/SBOX[10].sbox/U131  ( .A(n2601), .B(n2550), .Z(shift_row_out[18]) );
  XOR \b/SBOX[10].sbox/U130  ( .A(\b/SBOX[10].sbox/z[11] ), .B(n2604), .Z(
        n2550) );
  XOR \b/SBOX[10].sbox/U129  ( .A(n2552), .B(n2551), .Z(shift_row_out[19]) );
  XOR \b/SBOX[10].sbox/U128  ( .A(n2603), .B(n2553), .Z(n2551) );
  XOR \b/SBOX[10].sbox/U127  ( .A(\b/SBOX[10].sbox/z[5] ), .B(
        \b/SBOX[10].sbox/z[9] ), .Z(n2552) );
  XOR \b/SBOX[10].sbox/U126  ( .A(\b/SBOX[10].sbox/z[1] ), .B(
        \b/SBOX[10].sbox/z[2] ), .Z(n2553) );
  XOR \b/SBOX[10].sbox/U125  ( .A(n2602), .B(n2554), .Z(shift_row_out[20]) );
  XOR \b/SBOX[10].sbox/U124  ( .A(\b/SBOX[10].sbox/z[3] ), .B(n2603), .Z(n2554) );
  XOR \b/SBOX[10].sbox/U123  ( .A(n2604), .B(n2555), .Z(shift_row_out[23]) );
  XOR \b/SBOX[10].sbox/U122  ( .A(\b/SBOX[10].sbox/z[6] ), .B(
        \b/SBOX[10].sbox/z[9] ), .Z(n2555) );
  XOR \b/SBOX[10].sbox/U121  ( .A(n2557), .B(n2556), .Z(n2605) );
  XOR \b/SBOX[10].sbox/U120  ( .A(n2559), .B(n2558), .Z(n2556) );
  XOR \b/SBOX[10].sbox/U119  ( .A(msg[85]), .B(msg[81]), .Z(n2557) );
  XOR \b/SBOX[10].sbox/U118  ( .A(\b/SBOX[10].sbox/t[36] ), .B(
        \b/SBOX[10].sbox/t[39] ), .Z(n2558) );
  XOR \b/SBOX[10].sbox/U117  ( .A(\b/SBOX[10].sbox/t[3] ), .B(
        \b/SBOX[10].sbox/t[8] ), .Z(n2559) );
  XOR \b/SBOX[10].sbox/U116  ( .A(n2561), .B(n2560), .Z(
        \b/SBOX[10].sbox/t[41] ) );
  XOR \b/SBOX[10].sbox/U115  ( .A(n2605), .B(n2562), .Z(n2560) );
  XOR \b/SBOX[10].sbox/U114  ( .A(\b/SBOX[10].sbox/t[32] ), .B(msg[87]), .Z(
        n2561) );
  XOR \b/SBOX[10].sbox/U113  ( .A(\b/SBOX[10].sbox/t[5] ), .B(
        \b/SBOX[10].sbox/t[10] ), .Z(n2562) );
  XOR \b/SBOX[10].sbox/U112  ( .A(\b/SBOX[10].sbox/t[2] ), .B(msg[86]), .Z(
        n2606) );
  XOR \b/SBOX[10].sbox/U111  ( .A(n2564), .B(n2563), .Z(
        \b/SBOX[10].sbox/t[45] ) );
  XOR \b/SBOX[10].sbox/U110  ( .A(n2606), .B(n2565), .Z(n2563) );
  XOR \b/SBOX[10].sbox/U109  ( .A(msg[84]), .B(n2605), .Z(n2564) );
  XOR \b/SBOX[10].sbox/U108  ( .A(\b/SBOX[10].sbox/t[7] ), .B(
        \b/SBOX[10].sbox/t[28] ), .Z(n2565) );
  XOR \b/SBOX[10].sbox/U107  ( .A(n2606), .B(n2566), .Z(n2611) );
  XOR \b/SBOX[10].sbox/U106  ( .A(\b/SBOX[10].sbox/t[5] ), .B(msg[84]), .Z(
        n2566) );
  XOR \b/SBOX[10].sbox/U105  ( .A(msg[87]), .B(n2567), .Z(n2607) );
  XOR \b/SBOX[10].sbox/U104  ( .A(\b/SBOX[10].sbox/t[7] ), .B(
        \b/SBOX[10].sbox/t[10] ), .Z(n2567) );
  XOR \b/SBOX[10].sbox/U103  ( .A(n2569), .B(n2568), .Z(
        \b/SBOX[10].sbox/t[42] ) );
  XOR \b/SBOX[10].sbox/U102  ( .A(n2611), .B(n2607), .Z(n2568) );
  XOR \b/SBOX[10].sbox/U101  ( .A(\b/SBOX[10].sbox/t[28] ), .B(
        \b/SBOX[10].sbox/t[32] ), .Z(n2569) );
  XOR \b/SBOX[10].sbox/U100  ( .A(msg[81]), .B(n2570), .Z(n2609) );
  XOR \b/SBOX[10].sbox/U99  ( .A(msg[83]), .B(msg[82]), .Z(n2570) );
  XOR \b/SBOX[10].sbox/U98  ( .A(msg[85]), .B(n2609), .Z(
        \b/SBOX[10].sbox/y[16] ) );
  XOR \b/SBOX[10].sbox/U97  ( .A(\b/SBOX[10].sbox/y[16] ), .B(n2571), .Z(n2610) );
  XOR \b/SBOX[10].sbox/U96  ( .A(\b/SBOX[10].sbox/t[12] ), .B(
        \b/SBOX[10].sbox/t[15] ), .Z(n2571) );
  XOR \b/SBOX[10].sbox/U95  ( .A(n2610), .B(n2572), .Z(\b/SBOX[10].sbox/t[29] ) );
  XOR \b/SBOX[10].sbox/U94  ( .A(\b/SBOX[10].sbox/t[28] ), .B(n2611), .Z(n2572) );
  XOR \b/SBOX[10].sbox/U93  ( .A(msg[80]), .B(n2573), .Z(
        \b/SBOX[10].sbox/y[1] ) );
  XOR \b/SBOX[10].sbox/U92  ( .A(msg[86]), .B(msg[85]), .Z(n2573) );
  XOR \b/SBOX[10].sbox/U91  ( .A(msg[87]), .B(\b/SBOX[10].sbox/y[1] ), .Z(
        \b/SBOX[10].sbox/y[2] ) );
  XOR \b/SBOX[10].sbox/U90  ( .A(n2575), .B(n2574), .Z(\b/SBOX[10].sbox/t[25] ) );
  XOR \b/SBOX[10].sbox/U89  ( .A(n2577), .B(n2576), .Z(n2574) );
  XOR \b/SBOX[10].sbox/U88  ( .A(msg[87]), .B(msg[85]), .Z(n2575) );
  XOR \b/SBOX[10].sbox/U87  ( .A(\b/SBOX[10].sbox/t[13] ), .B(
        \b/SBOX[10].sbox/t[15] ), .Z(n2576) );
  XOR \b/SBOX[10].sbox/U86  ( .A(\b/SBOX[10].sbox/t[3] ), .B(
        \b/SBOX[10].sbox/t[5] ), .Z(n2577) );
  XOR \b/SBOX[10].sbox/U85  ( .A(\b/SBOX[10].sbox/t[39] ), .B(
        \b/SBOX[10].sbox/t[25] ), .Z(\b/SBOX[10].sbox/t[40] ) );
  XOR \b/SBOX[10].sbox/U84  ( .A(msg[81]), .B(\b/SBOX[10].sbox/y[1] ), .Z(
        \b/SBOX[10].sbox/y[5] ) );
  XOR \b/SBOX[10].sbox/U83  ( .A(n2579), .B(n2578), .Z(\b/SBOX[10].sbox/y[15] ) );
  XOR \b/SBOX[10].sbox/U82  ( .A(msg[83]), .B(msg[81]), .Z(n2578) );
  XOR \b/SBOX[10].sbox/U81  ( .A(msg[87]), .B(msg[84]), .Z(n2579) );
  XOR \b/SBOX[10].sbox/U80  ( .A(n2581), .B(n2580), .Z(\b/SBOX[10].sbox/t[21] ) );
  XOR \b/SBOX[10].sbox/U79  ( .A(n2583), .B(n2582), .Z(n2580) );
  XOR \b/SBOX[10].sbox/U78  ( .A(\b/SBOX[10].sbox/y[15] ), .B(n2606), .Z(n2581) );
  XOR \b/SBOX[10].sbox/U77  ( .A(\b/SBOX[10].sbox/t[13] ), .B(msg[82]), .Z(
        n2582) );
  XOR \b/SBOX[10].sbox/U76  ( .A(\b/SBOX[10].sbox/t[3] ), .B(
        \b/SBOX[10].sbox/t[12] ), .Z(n2583) );
  XOR \b/SBOX[10].sbox/U75  ( .A(\b/SBOX[10].sbox/t[21] ), .B(n2584), .Z(
        \b/SBOX[10].sbox/t[43] ) );
  XOR \b/SBOX[10].sbox/U74  ( .A(\b/SBOX[10].sbox/t[28] ), .B(
        \b/SBOX[10].sbox/t[39] ), .Z(n2584) );
  XOR \b/SBOX[10].sbox/U73  ( .A(n2610), .B(n2607), .Z(\b/SBOX[10].sbox/t[24] ) );
  XOR \b/SBOX[10].sbox/U72  ( .A(\b/SBOX[10].sbox/t[32] ), .B(
        \b/SBOX[10].sbox/t[24] ), .Z(\b/SBOX[10].sbox/t[33] ) );
  XOR \b/SBOX[10].sbox/U71  ( .A(msg[84]), .B(\b/SBOX[10].sbox/y[1] ), .Z(
        \b/SBOX[10].sbox/y[4] ) );
  XOR \b/SBOX[10].sbox/U70  ( .A(n2586), .B(n2585), .Z(\b/SBOX[10].sbox/t[30] ) );
  XOR \b/SBOX[10].sbox/U69  ( .A(msg[81]), .B(n2587), .Z(n2585) );
  XOR \b/SBOX[10].sbox/U68  ( .A(\b/SBOX[10].sbox/t[13] ), .B(
        \b/SBOX[10].sbox/t[15] ), .Z(n2586) );
  XOR \b/SBOX[10].sbox/U67  ( .A(\b/SBOX[10].sbox/t[8] ), .B(
        \b/SBOX[10].sbox/t[10] ), .Z(n2587) );
  XOR \b/SBOX[10].sbox/U66  ( .A(\b/SBOX[10].sbox/t[30] ), .B(n2588), .Z(
        \b/SBOX[10].sbox/t[37] ) );
  XOR \b/SBOX[10].sbox/U65  ( .A(\b/SBOX[10].sbox/t[32] ), .B(
        \b/SBOX[10].sbox/t[36] ), .Z(n2588) );
  XOR \b/SBOX[10].sbox/U64  ( .A(msg[87]), .B(msg[82]), .Z(n2608) );
  XOR \b/SBOX[10].sbox/U63  ( .A(\b/SBOX[10].sbox/y[5] ), .B(n2608), .Z(
        \b/SBOX[10].sbox/y[3] ) );
  XOR \b/SBOX[10].sbox/U62  ( .A(n2590), .B(n2589), .Z(\b/SBOX[10].sbox/t[23] ) );
  XOR \b/SBOX[10].sbox/U61  ( .A(n2592), .B(n2591), .Z(n2589) );
  XOR \b/SBOX[10].sbox/U60  ( .A(n2608), .B(n2593), .Z(n2590) );
  XOR \b/SBOX[10].sbox/U59  ( .A(msg[85]), .B(msg[83]), .Z(n2591) );
  XOR \b/SBOX[10].sbox/U58  ( .A(\b/SBOX[10].sbox/t[12] ), .B(
        \b/SBOX[10].sbox/t[13] ), .Z(n2592) );
  XOR \b/SBOX[10].sbox/U57  ( .A(\b/SBOX[10].sbox/t[7] ), .B(
        \b/SBOX[10].sbox/t[8] ), .Z(n2593) );
  XOR \b/SBOX[10].sbox/U56  ( .A(\b/SBOX[10].sbox/t[36] ), .B(
        \b/SBOX[10].sbox/t[23] ), .Z(\b/SBOX[10].sbox/t[44] ) );
  XOR \b/SBOX[10].sbox/U55  ( .A(n2608), .B(n2594), .Z(\b/SBOX[10].sbox/y[12] ) );
  XOR \b/SBOX[10].sbox/U54  ( .A(msg[84]), .B(msg[81]), .Z(n2594) );
  XOR \b/SBOX[10].sbox/U53  ( .A(\b/SBOX[10].sbox/y[15] ), .B(n2595), .Z(
        \b/SBOX[10].sbox/y[10] ) );
  XOR \b/SBOX[10].sbox/U52  ( .A(msg[86]), .B(msg[85]), .Z(n2595) );
  XOR \b/SBOX[10].sbox/U51  ( .A(n2608), .B(n2596), .Z(\b/SBOX[10].sbox/y[17] ) );
  XOR \b/SBOX[10].sbox/U50  ( .A(msg[85]), .B(msg[84]), .Z(n2596) );
  XOR \b/SBOX[10].sbox/U49  ( .A(msg[86]), .B(n2609), .Z(
        \b/SBOX[10].sbox/y[11] ) );
  XOR \b/SBOX[10].sbox/U48  ( .A(msg[80]), .B(\b/SBOX[10].sbox/y[11] ), .Z(
        \b/SBOX[10].sbox/y[7] ) );
  XOR \b/SBOX[10].sbox/U47  ( .A(msg[80]), .B(\b/SBOX[10].sbox/y[15] ), .Z(
        \b/SBOX[10].sbox/y[6] ) );
  XOR \b/SBOX[10].sbox/U46  ( .A(\b/SBOX[10].sbox/t[26] ), .B(
        \b/SBOX[10].sbox/t[24] ), .Z(\b/SBOX[10].sbox/t[27] ) );
  XOR \b/SBOX[10].sbox/U45  ( .A(\b/SBOX[10].sbox/t[36] ), .B(
        \b/SBOX[10].sbox/t[27] ), .Z(\b/SBOX[10].sbox/t[38] ) );
  XOR \b/SBOX[10].sbox/U44  ( .A(n2610), .B(n2597), .Z(\b/SBOX[10].sbox/t[31] ) );
  XOR \b/SBOX[10].sbox/U43  ( .A(\b/SBOX[10].sbox/t[26] ), .B(n2611), .Z(n2597) );
  XOR \b/SBOX[9].sbox/U157  ( .A(\b/SBOX[9].sbox/z[12] ), .B(n2454), .Z(n2518)
         );
  XOR \b/SBOX[9].sbox/U156  ( .A(\b/SBOX[9].sbox/z[0] ), .B(
        \b/SBOX[9].sbox/z[2] ), .Z(n2454) );
  XOR \b/SBOX[9].sbox/U155  ( .A(n2456), .B(n2455), .Z(n2517) );
  XOR \b/SBOX[9].sbox/U154  ( .A(\b/SBOX[9].sbox/z[15] ), .B(
        \b/SBOX[9].sbox/z[16] ), .Z(n2455) );
  XOR \b/SBOX[9].sbox/U153  ( .A(\b/SBOX[9].sbox/z[5] ), .B(
        \b/SBOX[9].sbox/z[13] ), .Z(n2456) );
  XOR \b/SBOX[9].sbox/U152  ( .A(n2517), .B(n2457), .Z(n2531) );
  XOR \b/SBOX[9].sbox/U151  ( .A(\b/SBOX[9].sbox/z[3] ), .B(n2518), .Z(n2457)
         );
  XOR \b/SBOX[9].sbox/U150  ( .A(n2459), .B(n2458), .Z(n2532) );
  XOR \b/SBOX[9].sbox/U149  ( .A(n2517), .B(n2460), .Z(n2458) );
  XOR \b/SBOX[9].sbox/U148  ( .A(\b/SBOX[9].sbox/z[8] ), .B(
        \b/SBOX[9].sbox/z[12] ), .Z(n2459) );
  XOR \b/SBOX[9].sbox/U147  ( .A(\b/SBOX[9].sbox/z[4] ), .B(
        \b/SBOX[9].sbox/z[7] ), .Z(n2460) );
  XOR \b/SBOX[9].sbox/U146  ( .A(n2518), .B(n2461), .Z(n2520) );
  XOR \b/SBOX[9].sbox/U145  ( .A(\b/SBOX[9].sbox/z[8] ), .B(
        \b/SBOX[9].sbox/z[14] ), .Z(n2461) );
  XOR \b/SBOX[9].sbox/U144  ( .A(n2463), .B(n2462), .Z(n2533) );
  XOR \b/SBOX[9].sbox/U143  ( .A(\b/SBOX[9].sbox/z[17] ), .B(n2520), .Z(n2462)
         );
  XOR \b/SBOX[9].sbox/U142  ( .A(\b/SBOX[9].sbox/z[6] ), .B(
        \b/SBOX[9].sbox/z[15] ), .Z(n2463) );
  XOR \b/SBOX[9].sbox/U141  ( .A(\b/SBOX[9].sbox/z[9] ), .B(n2464), .Z(n2521)
         );
  XOR \b/SBOX[9].sbox/U140  ( .A(\b/SBOX[9].sbox/z[0] ), .B(
        \b/SBOX[9].sbox/z[1] ), .Z(n2464) );
  XOR \b/SBOX[9].sbox/U139  ( .A(\b/SBOX[9].sbox/z[16] ), .B(n2465), .Z(n2519)
         );
  XOR \b/SBOX[9].sbox/U138  ( .A(\b/SBOX[9].sbox/z[10] ), .B(
        \b/SBOX[9].sbox/z[15] ), .Z(n2465) );
  XOR \b/SBOX[9].sbox/U137  ( .A(n2467), .B(n2466), .Z(n2534) );
  XOR \b/SBOX[9].sbox/U136  ( .A(n2521), .B(n2519), .Z(n2466) );
  XOR \b/SBOX[9].sbox/U135  ( .A(\b/SBOX[9].sbox/z[6] ), .B(
        \b/SBOX[9].sbox/z[7] ), .Z(n2467) );
  XOR \b/SBOX[9].sbox/U134  ( .A(\b/SBOX[9].sbox/z[4] ), .B(n2519), .Z(n2522)
         );
  XOR \b/SBOX[9].sbox/U133  ( .A(n2522), .B(n2468), .Z(n2523) );
  XOR \b/SBOX[9].sbox/U132  ( .A(\b/SBOX[9].sbox/z[3] ), .B(
        \b/SBOX[9].sbox/z[7] ), .Z(n2468) );
  XOR \b/SBOX[9].sbox/U131  ( .A(n2520), .B(n2469), .Z(shift_row_out[42]) );
  XOR \b/SBOX[9].sbox/U130  ( .A(\b/SBOX[9].sbox/z[11] ), .B(n2523), .Z(n2469)
         );
  XOR \b/SBOX[9].sbox/U129  ( .A(n2471), .B(n2470), .Z(shift_row_out[43]) );
  XOR \b/SBOX[9].sbox/U128  ( .A(n2522), .B(n2472), .Z(n2470) );
  XOR \b/SBOX[9].sbox/U127  ( .A(\b/SBOX[9].sbox/z[5] ), .B(
        \b/SBOX[9].sbox/z[9] ), .Z(n2471) );
  XOR \b/SBOX[9].sbox/U126  ( .A(\b/SBOX[9].sbox/z[1] ), .B(
        \b/SBOX[9].sbox/z[2] ), .Z(n2472) );
  XOR \b/SBOX[9].sbox/U125  ( .A(n2521), .B(n2473), .Z(shift_row_out[44]) );
  XOR \b/SBOX[9].sbox/U124  ( .A(\b/SBOX[9].sbox/z[3] ), .B(n2522), .Z(n2473)
         );
  XOR \b/SBOX[9].sbox/U123  ( .A(n2523), .B(n2474), .Z(shift_row_out[47]) );
  XOR \b/SBOX[9].sbox/U122  ( .A(\b/SBOX[9].sbox/z[6] ), .B(
        \b/SBOX[9].sbox/z[9] ), .Z(n2474) );
  XOR \b/SBOX[9].sbox/U121  ( .A(n2476), .B(n2475), .Z(n2524) );
  XOR \b/SBOX[9].sbox/U120  ( .A(n2478), .B(n2477), .Z(n2475) );
  XOR \b/SBOX[9].sbox/U119  ( .A(msg[77]), .B(msg[73]), .Z(n2476) );
  XOR \b/SBOX[9].sbox/U118  ( .A(\b/SBOX[9].sbox/t[36] ), .B(
        \b/SBOX[9].sbox/t[39] ), .Z(n2477) );
  XOR \b/SBOX[9].sbox/U117  ( .A(\b/SBOX[9].sbox/t[3] ), .B(
        \b/SBOX[9].sbox/t[8] ), .Z(n2478) );
  XOR \b/SBOX[9].sbox/U116  ( .A(n2480), .B(n2479), .Z(\b/SBOX[9].sbox/t[41] )
         );
  XOR \b/SBOX[9].sbox/U115  ( .A(n2524), .B(n2481), .Z(n2479) );
  XOR \b/SBOX[9].sbox/U114  ( .A(\b/SBOX[9].sbox/t[32] ), .B(msg[79]), .Z(
        n2480) );
  XOR \b/SBOX[9].sbox/U113  ( .A(\b/SBOX[9].sbox/t[5] ), .B(
        \b/SBOX[9].sbox/t[10] ), .Z(n2481) );
  XOR \b/SBOX[9].sbox/U112  ( .A(\b/SBOX[9].sbox/t[2] ), .B(msg[78]), .Z(n2525) );
  XOR \b/SBOX[9].sbox/U111  ( .A(n2483), .B(n2482), .Z(\b/SBOX[9].sbox/t[45] )
         );
  XOR \b/SBOX[9].sbox/U110  ( .A(n2525), .B(n2484), .Z(n2482) );
  XOR \b/SBOX[9].sbox/U109  ( .A(msg[76]), .B(n2524), .Z(n2483) );
  XOR \b/SBOX[9].sbox/U108  ( .A(\b/SBOX[9].sbox/t[7] ), .B(
        \b/SBOX[9].sbox/t[28] ), .Z(n2484) );
  XOR \b/SBOX[9].sbox/U107  ( .A(n2525), .B(n2485), .Z(n2530) );
  XOR \b/SBOX[9].sbox/U106  ( .A(\b/SBOX[9].sbox/t[5] ), .B(msg[76]), .Z(n2485) );
  XOR \b/SBOX[9].sbox/U105  ( .A(msg[79]), .B(n2486), .Z(n2526) );
  XOR \b/SBOX[9].sbox/U104  ( .A(\b/SBOX[9].sbox/t[7] ), .B(
        \b/SBOX[9].sbox/t[10] ), .Z(n2486) );
  XOR \b/SBOX[9].sbox/U103  ( .A(n2488), .B(n2487), .Z(\b/SBOX[9].sbox/t[42] )
         );
  XOR \b/SBOX[9].sbox/U102  ( .A(n2530), .B(n2526), .Z(n2487) );
  XOR \b/SBOX[9].sbox/U101  ( .A(\b/SBOX[9].sbox/t[28] ), .B(
        \b/SBOX[9].sbox/t[32] ), .Z(n2488) );
  XOR \b/SBOX[9].sbox/U100  ( .A(msg[73]), .B(n2489), .Z(n2528) );
  XOR \b/SBOX[9].sbox/U99  ( .A(msg[75]), .B(msg[74]), .Z(n2489) );
  XOR \b/SBOX[9].sbox/U98  ( .A(msg[77]), .B(n2528), .Z(\b/SBOX[9].sbox/y[16] ) );
  XOR \b/SBOX[9].sbox/U97  ( .A(\b/SBOX[9].sbox/y[16] ), .B(n2490), .Z(n2529)
         );
  XOR \b/SBOX[9].sbox/U96  ( .A(\b/SBOX[9].sbox/t[12] ), .B(
        \b/SBOX[9].sbox/t[15] ), .Z(n2490) );
  XOR \b/SBOX[9].sbox/U95  ( .A(n2529), .B(n2491), .Z(\b/SBOX[9].sbox/t[29] )
         );
  XOR \b/SBOX[9].sbox/U94  ( .A(\b/SBOX[9].sbox/t[28] ), .B(n2530), .Z(n2491)
         );
  XOR \b/SBOX[9].sbox/U93  ( .A(msg[72]), .B(n2492), .Z(\b/SBOX[9].sbox/y[1] )
         );
  XOR \b/SBOX[9].sbox/U92  ( .A(msg[78]), .B(msg[77]), .Z(n2492) );
  XOR \b/SBOX[9].sbox/U91  ( .A(msg[79]), .B(\b/SBOX[9].sbox/y[1] ), .Z(
        \b/SBOX[9].sbox/y[2] ) );
  XOR \b/SBOX[9].sbox/U90  ( .A(n2494), .B(n2493), .Z(\b/SBOX[9].sbox/t[25] )
         );
  XOR \b/SBOX[9].sbox/U89  ( .A(n2496), .B(n2495), .Z(n2493) );
  XOR \b/SBOX[9].sbox/U88  ( .A(msg[79]), .B(msg[77]), .Z(n2494) );
  XOR \b/SBOX[9].sbox/U87  ( .A(\b/SBOX[9].sbox/t[13] ), .B(
        \b/SBOX[9].sbox/t[15] ), .Z(n2495) );
  XOR \b/SBOX[9].sbox/U86  ( .A(\b/SBOX[9].sbox/t[3] ), .B(
        \b/SBOX[9].sbox/t[5] ), .Z(n2496) );
  XOR \b/SBOX[9].sbox/U85  ( .A(\b/SBOX[9].sbox/t[39] ), .B(
        \b/SBOX[9].sbox/t[25] ), .Z(\b/SBOX[9].sbox/t[40] ) );
  XOR \b/SBOX[9].sbox/U84  ( .A(msg[73]), .B(\b/SBOX[9].sbox/y[1] ), .Z(
        \b/SBOX[9].sbox/y[5] ) );
  XOR \b/SBOX[9].sbox/U83  ( .A(n2498), .B(n2497), .Z(\b/SBOX[9].sbox/y[15] )
         );
  XOR \b/SBOX[9].sbox/U82  ( .A(msg[75]), .B(msg[73]), .Z(n2497) );
  XOR \b/SBOX[9].sbox/U81  ( .A(msg[79]), .B(msg[76]), .Z(n2498) );
  XOR \b/SBOX[9].sbox/U80  ( .A(n2500), .B(n2499), .Z(\b/SBOX[9].sbox/t[21] )
         );
  XOR \b/SBOX[9].sbox/U79  ( .A(n2502), .B(n2501), .Z(n2499) );
  XOR \b/SBOX[9].sbox/U78  ( .A(\b/SBOX[9].sbox/y[15] ), .B(n2525), .Z(n2500)
         );
  XOR \b/SBOX[9].sbox/U77  ( .A(\b/SBOX[9].sbox/t[13] ), .B(msg[74]), .Z(n2501) );
  XOR \b/SBOX[9].sbox/U76  ( .A(\b/SBOX[9].sbox/t[3] ), .B(
        \b/SBOX[9].sbox/t[12] ), .Z(n2502) );
  XOR \b/SBOX[9].sbox/U75  ( .A(\b/SBOX[9].sbox/t[21] ), .B(n2503), .Z(
        \b/SBOX[9].sbox/t[43] ) );
  XOR \b/SBOX[9].sbox/U74  ( .A(\b/SBOX[9].sbox/t[28] ), .B(
        \b/SBOX[9].sbox/t[39] ), .Z(n2503) );
  XOR \b/SBOX[9].sbox/U73  ( .A(n2529), .B(n2526), .Z(\b/SBOX[9].sbox/t[24] )
         );
  XOR \b/SBOX[9].sbox/U72  ( .A(\b/SBOX[9].sbox/t[32] ), .B(
        \b/SBOX[9].sbox/t[24] ), .Z(\b/SBOX[9].sbox/t[33] ) );
  XOR \b/SBOX[9].sbox/U71  ( .A(msg[76]), .B(\b/SBOX[9].sbox/y[1] ), .Z(
        \b/SBOX[9].sbox/y[4] ) );
  XOR \b/SBOX[9].sbox/U70  ( .A(n2505), .B(n2504), .Z(\b/SBOX[9].sbox/t[30] )
         );
  XOR \b/SBOX[9].sbox/U69  ( .A(msg[73]), .B(n2506), .Z(n2504) );
  XOR \b/SBOX[9].sbox/U68  ( .A(\b/SBOX[9].sbox/t[13] ), .B(
        \b/SBOX[9].sbox/t[15] ), .Z(n2505) );
  XOR \b/SBOX[9].sbox/U67  ( .A(\b/SBOX[9].sbox/t[8] ), .B(
        \b/SBOX[9].sbox/t[10] ), .Z(n2506) );
  XOR \b/SBOX[9].sbox/U66  ( .A(\b/SBOX[9].sbox/t[30] ), .B(n2507), .Z(
        \b/SBOX[9].sbox/t[37] ) );
  XOR \b/SBOX[9].sbox/U65  ( .A(\b/SBOX[9].sbox/t[32] ), .B(
        \b/SBOX[9].sbox/t[36] ), .Z(n2507) );
  XOR \b/SBOX[9].sbox/U64  ( .A(msg[79]), .B(msg[74]), .Z(n2527) );
  XOR \b/SBOX[9].sbox/U63  ( .A(\b/SBOX[9].sbox/y[5] ), .B(n2527), .Z(
        \b/SBOX[9].sbox/y[3] ) );
  XOR \b/SBOX[9].sbox/U62  ( .A(n2509), .B(n2508), .Z(\b/SBOX[9].sbox/t[23] )
         );
  XOR \b/SBOX[9].sbox/U61  ( .A(n2511), .B(n2510), .Z(n2508) );
  XOR \b/SBOX[9].sbox/U60  ( .A(n2527), .B(n2512), .Z(n2509) );
  XOR \b/SBOX[9].sbox/U59  ( .A(msg[77]), .B(msg[75]), .Z(n2510) );
  XOR \b/SBOX[9].sbox/U58  ( .A(\b/SBOX[9].sbox/t[12] ), .B(
        \b/SBOX[9].sbox/t[13] ), .Z(n2511) );
  XOR \b/SBOX[9].sbox/U57  ( .A(\b/SBOX[9].sbox/t[7] ), .B(
        \b/SBOX[9].sbox/t[8] ), .Z(n2512) );
  XOR \b/SBOX[9].sbox/U56  ( .A(\b/SBOX[9].sbox/t[36] ), .B(
        \b/SBOX[9].sbox/t[23] ), .Z(\b/SBOX[9].sbox/t[44] ) );
  XOR \b/SBOX[9].sbox/U55  ( .A(n2527), .B(n2513), .Z(\b/SBOX[9].sbox/y[12] )
         );
  XOR \b/SBOX[9].sbox/U54  ( .A(msg[76]), .B(msg[73]), .Z(n2513) );
  XOR \b/SBOX[9].sbox/U53  ( .A(\b/SBOX[9].sbox/y[15] ), .B(n2514), .Z(
        \b/SBOX[9].sbox/y[10] ) );
  XOR \b/SBOX[9].sbox/U52  ( .A(msg[78]), .B(msg[77]), .Z(n2514) );
  XOR \b/SBOX[9].sbox/U51  ( .A(n2527), .B(n2515), .Z(\b/SBOX[9].sbox/y[17] )
         );
  XOR \b/SBOX[9].sbox/U50  ( .A(msg[77]), .B(msg[76]), .Z(n2515) );
  XOR \b/SBOX[9].sbox/U49  ( .A(msg[78]), .B(n2528), .Z(\b/SBOX[9].sbox/y[11] ) );
  XOR \b/SBOX[9].sbox/U48  ( .A(msg[72]), .B(\b/SBOX[9].sbox/y[11] ), .Z(
        \b/SBOX[9].sbox/y[7] ) );
  XOR \b/SBOX[9].sbox/U47  ( .A(msg[72]), .B(\b/SBOX[9].sbox/y[15] ), .Z(
        \b/SBOX[9].sbox/y[6] ) );
  XOR \b/SBOX[9].sbox/U46  ( .A(\b/SBOX[9].sbox/t[26] ), .B(
        \b/SBOX[9].sbox/t[24] ), .Z(\b/SBOX[9].sbox/t[27] ) );
  XOR \b/SBOX[9].sbox/U45  ( .A(\b/SBOX[9].sbox/t[36] ), .B(
        \b/SBOX[9].sbox/t[27] ), .Z(\b/SBOX[9].sbox/t[38] ) );
  XOR \b/SBOX[9].sbox/U44  ( .A(n2529), .B(n2516), .Z(\b/SBOX[9].sbox/t[31] )
         );
  XOR \b/SBOX[9].sbox/U43  ( .A(\b/SBOX[9].sbox/t[26] ), .B(n2530), .Z(n2516)
         );
  XOR \b/SBOX[8].sbox/U157  ( .A(\b/SBOX[8].sbox/z[12] ), .B(n2373), .Z(n2437)
         );
  XOR \b/SBOX[8].sbox/U156  ( .A(\b/SBOX[8].sbox/z[0] ), .B(
        \b/SBOX[8].sbox/z[2] ), .Z(n2373) );
  XOR \b/SBOX[8].sbox/U155  ( .A(n2375), .B(n2374), .Z(n2436) );
  XOR \b/SBOX[8].sbox/U154  ( .A(\b/SBOX[8].sbox/z[15] ), .B(
        \b/SBOX[8].sbox/z[16] ), .Z(n2374) );
  XOR \b/SBOX[8].sbox/U153  ( .A(\b/SBOX[8].sbox/z[5] ), .B(
        \b/SBOX[8].sbox/z[13] ), .Z(n2375) );
  XOR \b/SBOX[8].sbox/U152  ( .A(n2436), .B(n2376), .Z(n2450) );
  XOR \b/SBOX[8].sbox/U151  ( .A(\b/SBOX[8].sbox/z[3] ), .B(n2437), .Z(n2376)
         );
  XOR \b/SBOX[8].sbox/U150  ( .A(n2378), .B(n2377), .Z(n2451) );
  XOR \b/SBOX[8].sbox/U149  ( .A(n2436), .B(n2379), .Z(n2377) );
  XOR \b/SBOX[8].sbox/U148  ( .A(\b/SBOX[8].sbox/z[8] ), .B(
        \b/SBOX[8].sbox/z[12] ), .Z(n2378) );
  XOR \b/SBOX[8].sbox/U147  ( .A(\b/SBOX[8].sbox/z[4] ), .B(
        \b/SBOX[8].sbox/z[7] ), .Z(n2379) );
  XOR \b/SBOX[8].sbox/U146  ( .A(n2437), .B(n2380), .Z(n2439) );
  XOR \b/SBOX[8].sbox/U145  ( .A(\b/SBOX[8].sbox/z[8] ), .B(
        \b/SBOX[8].sbox/z[14] ), .Z(n2380) );
  XOR \b/SBOX[8].sbox/U144  ( .A(n2382), .B(n2381), .Z(n2452) );
  XOR \b/SBOX[8].sbox/U143  ( .A(\b/SBOX[8].sbox/z[17] ), .B(n2439), .Z(n2381)
         );
  XOR \b/SBOX[8].sbox/U142  ( .A(\b/SBOX[8].sbox/z[6] ), .B(
        \b/SBOX[8].sbox/z[15] ), .Z(n2382) );
  XOR \b/SBOX[8].sbox/U141  ( .A(\b/SBOX[8].sbox/z[9] ), .B(n2383), .Z(n2440)
         );
  XOR \b/SBOX[8].sbox/U140  ( .A(\b/SBOX[8].sbox/z[0] ), .B(
        \b/SBOX[8].sbox/z[1] ), .Z(n2383) );
  XOR \b/SBOX[8].sbox/U139  ( .A(\b/SBOX[8].sbox/z[16] ), .B(n2384), .Z(n2438)
         );
  XOR \b/SBOX[8].sbox/U138  ( .A(\b/SBOX[8].sbox/z[10] ), .B(
        \b/SBOX[8].sbox/z[15] ), .Z(n2384) );
  XOR \b/SBOX[8].sbox/U137  ( .A(n2386), .B(n2385), .Z(n2453) );
  XOR \b/SBOX[8].sbox/U136  ( .A(n2440), .B(n2438), .Z(n2385) );
  XOR \b/SBOX[8].sbox/U135  ( .A(\b/SBOX[8].sbox/z[6] ), .B(
        \b/SBOX[8].sbox/z[7] ), .Z(n2386) );
  XOR \b/SBOX[8].sbox/U134  ( .A(\b/SBOX[8].sbox/z[4] ), .B(n2438), .Z(n2441)
         );
  XOR \b/SBOX[8].sbox/U133  ( .A(n2441), .B(n2387), .Z(n2442) );
  XOR \b/SBOX[8].sbox/U132  ( .A(\b/SBOX[8].sbox/z[3] ), .B(
        \b/SBOX[8].sbox/z[7] ), .Z(n2387) );
  XOR \b/SBOX[8].sbox/U131  ( .A(n2439), .B(n2388), .Z(shift_row_out[66]) );
  XOR \b/SBOX[8].sbox/U130  ( .A(\b/SBOX[8].sbox/z[11] ), .B(n2442), .Z(n2388)
         );
  XOR \b/SBOX[8].sbox/U129  ( .A(n2390), .B(n2389), .Z(shift_row_out[67]) );
  XOR \b/SBOX[8].sbox/U128  ( .A(n2441), .B(n2391), .Z(n2389) );
  XOR \b/SBOX[8].sbox/U127  ( .A(\b/SBOX[8].sbox/z[5] ), .B(
        \b/SBOX[8].sbox/z[9] ), .Z(n2390) );
  XOR \b/SBOX[8].sbox/U126  ( .A(\b/SBOX[8].sbox/z[1] ), .B(
        \b/SBOX[8].sbox/z[2] ), .Z(n2391) );
  XOR \b/SBOX[8].sbox/U125  ( .A(n2440), .B(n2392), .Z(shift_row_out[68]) );
  XOR \b/SBOX[8].sbox/U124  ( .A(\b/SBOX[8].sbox/z[3] ), .B(n2441), .Z(n2392)
         );
  XOR \b/SBOX[8].sbox/U123  ( .A(n2442), .B(n2393), .Z(shift_row_out[71]) );
  XOR \b/SBOX[8].sbox/U122  ( .A(\b/SBOX[8].sbox/z[6] ), .B(
        \b/SBOX[8].sbox/z[9] ), .Z(n2393) );
  XOR \b/SBOX[8].sbox/U121  ( .A(n2395), .B(n2394), .Z(n2443) );
  XOR \b/SBOX[8].sbox/U120  ( .A(n2397), .B(n2396), .Z(n2394) );
  XOR \b/SBOX[8].sbox/U119  ( .A(msg[69]), .B(msg[65]), .Z(n2395) );
  XOR \b/SBOX[8].sbox/U118  ( .A(\b/SBOX[8].sbox/t[36] ), .B(
        \b/SBOX[8].sbox/t[39] ), .Z(n2396) );
  XOR \b/SBOX[8].sbox/U117  ( .A(\b/SBOX[8].sbox/t[3] ), .B(
        \b/SBOX[8].sbox/t[8] ), .Z(n2397) );
  XOR \b/SBOX[8].sbox/U116  ( .A(n2399), .B(n2398), .Z(\b/SBOX[8].sbox/t[41] )
         );
  XOR \b/SBOX[8].sbox/U115  ( .A(n2443), .B(n2400), .Z(n2398) );
  XOR \b/SBOX[8].sbox/U114  ( .A(\b/SBOX[8].sbox/t[32] ), .B(msg[71]), .Z(
        n2399) );
  XOR \b/SBOX[8].sbox/U113  ( .A(\b/SBOX[8].sbox/t[5] ), .B(
        \b/SBOX[8].sbox/t[10] ), .Z(n2400) );
  XOR \b/SBOX[8].sbox/U112  ( .A(\b/SBOX[8].sbox/t[2] ), .B(msg[70]), .Z(n2444) );
  XOR \b/SBOX[8].sbox/U111  ( .A(n2402), .B(n2401), .Z(\b/SBOX[8].sbox/t[45] )
         );
  XOR \b/SBOX[8].sbox/U110  ( .A(n2444), .B(n2403), .Z(n2401) );
  XOR \b/SBOX[8].sbox/U109  ( .A(msg[68]), .B(n2443), .Z(n2402) );
  XOR \b/SBOX[8].sbox/U108  ( .A(\b/SBOX[8].sbox/t[7] ), .B(
        \b/SBOX[8].sbox/t[28] ), .Z(n2403) );
  XOR \b/SBOX[8].sbox/U107  ( .A(n2444), .B(n2404), .Z(n2449) );
  XOR \b/SBOX[8].sbox/U106  ( .A(\b/SBOX[8].sbox/t[5] ), .B(msg[68]), .Z(n2404) );
  XOR \b/SBOX[8].sbox/U105  ( .A(msg[71]), .B(n2405), .Z(n2445) );
  XOR \b/SBOX[8].sbox/U104  ( .A(\b/SBOX[8].sbox/t[7] ), .B(
        \b/SBOX[8].sbox/t[10] ), .Z(n2405) );
  XOR \b/SBOX[8].sbox/U103  ( .A(n2407), .B(n2406), .Z(\b/SBOX[8].sbox/t[42] )
         );
  XOR \b/SBOX[8].sbox/U102  ( .A(n2449), .B(n2445), .Z(n2406) );
  XOR \b/SBOX[8].sbox/U101  ( .A(\b/SBOX[8].sbox/t[28] ), .B(
        \b/SBOX[8].sbox/t[32] ), .Z(n2407) );
  XOR \b/SBOX[8].sbox/U100  ( .A(msg[65]), .B(n2408), .Z(n2447) );
  XOR \b/SBOX[8].sbox/U99  ( .A(msg[67]), .B(msg[66]), .Z(n2408) );
  XOR \b/SBOX[8].sbox/U98  ( .A(msg[69]), .B(n2447), .Z(\b/SBOX[8].sbox/y[16] ) );
  XOR \b/SBOX[8].sbox/U97  ( .A(\b/SBOX[8].sbox/y[16] ), .B(n2409), .Z(n2448)
         );
  XOR \b/SBOX[8].sbox/U96  ( .A(\b/SBOX[8].sbox/t[12] ), .B(
        \b/SBOX[8].sbox/t[15] ), .Z(n2409) );
  XOR \b/SBOX[8].sbox/U95  ( .A(n2448), .B(n2410), .Z(\b/SBOX[8].sbox/t[29] )
         );
  XOR \b/SBOX[8].sbox/U94  ( .A(\b/SBOX[8].sbox/t[28] ), .B(n2449), .Z(n2410)
         );
  XOR \b/SBOX[8].sbox/U93  ( .A(msg[64]), .B(n2411), .Z(\b/SBOX[8].sbox/y[1] )
         );
  XOR \b/SBOX[8].sbox/U92  ( .A(msg[70]), .B(msg[69]), .Z(n2411) );
  XOR \b/SBOX[8].sbox/U91  ( .A(msg[71]), .B(\b/SBOX[8].sbox/y[1] ), .Z(
        \b/SBOX[8].sbox/y[2] ) );
  XOR \b/SBOX[8].sbox/U90  ( .A(n2413), .B(n2412), .Z(\b/SBOX[8].sbox/t[25] )
         );
  XOR \b/SBOX[8].sbox/U89  ( .A(n2415), .B(n2414), .Z(n2412) );
  XOR \b/SBOX[8].sbox/U88  ( .A(msg[71]), .B(msg[69]), .Z(n2413) );
  XOR \b/SBOX[8].sbox/U87  ( .A(\b/SBOX[8].sbox/t[13] ), .B(
        \b/SBOX[8].sbox/t[15] ), .Z(n2414) );
  XOR \b/SBOX[8].sbox/U86  ( .A(\b/SBOX[8].sbox/t[3] ), .B(
        \b/SBOX[8].sbox/t[5] ), .Z(n2415) );
  XOR \b/SBOX[8].sbox/U85  ( .A(\b/SBOX[8].sbox/t[39] ), .B(
        \b/SBOX[8].sbox/t[25] ), .Z(\b/SBOX[8].sbox/t[40] ) );
  XOR \b/SBOX[8].sbox/U84  ( .A(msg[65]), .B(\b/SBOX[8].sbox/y[1] ), .Z(
        \b/SBOX[8].sbox/y[5] ) );
  XOR \b/SBOX[8].sbox/U83  ( .A(n2417), .B(n2416), .Z(\b/SBOX[8].sbox/y[15] )
         );
  XOR \b/SBOX[8].sbox/U82  ( .A(msg[67]), .B(msg[65]), .Z(n2416) );
  XOR \b/SBOX[8].sbox/U81  ( .A(msg[71]), .B(msg[68]), .Z(n2417) );
  XOR \b/SBOX[8].sbox/U80  ( .A(n2419), .B(n2418), .Z(\b/SBOX[8].sbox/t[21] )
         );
  XOR \b/SBOX[8].sbox/U79  ( .A(n2421), .B(n2420), .Z(n2418) );
  XOR \b/SBOX[8].sbox/U78  ( .A(\b/SBOX[8].sbox/y[15] ), .B(n2444), .Z(n2419)
         );
  XOR \b/SBOX[8].sbox/U77  ( .A(\b/SBOX[8].sbox/t[13] ), .B(msg[66]), .Z(n2420) );
  XOR \b/SBOX[8].sbox/U76  ( .A(\b/SBOX[8].sbox/t[3] ), .B(
        \b/SBOX[8].sbox/t[12] ), .Z(n2421) );
  XOR \b/SBOX[8].sbox/U75  ( .A(\b/SBOX[8].sbox/t[21] ), .B(n2422), .Z(
        \b/SBOX[8].sbox/t[43] ) );
  XOR \b/SBOX[8].sbox/U74  ( .A(\b/SBOX[8].sbox/t[28] ), .B(
        \b/SBOX[8].sbox/t[39] ), .Z(n2422) );
  XOR \b/SBOX[8].sbox/U73  ( .A(n2448), .B(n2445), .Z(\b/SBOX[8].sbox/t[24] )
         );
  XOR \b/SBOX[8].sbox/U72  ( .A(\b/SBOX[8].sbox/t[32] ), .B(
        \b/SBOX[8].sbox/t[24] ), .Z(\b/SBOX[8].sbox/t[33] ) );
  XOR \b/SBOX[8].sbox/U71  ( .A(msg[68]), .B(\b/SBOX[8].sbox/y[1] ), .Z(
        \b/SBOX[8].sbox/y[4] ) );
  XOR \b/SBOX[8].sbox/U70  ( .A(n2424), .B(n2423), .Z(\b/SBOX[8].sbox/t[30] )
         );
  XOR \b/SBOX[8].sbox/U69  ( .A(msg[65]), .B(n2425), .Z(n2423) );
  XOR \b/SBOX[8].sbox/U68  ( .A(\b/SBOX[8].sbox/t[13] ), .B(
        \b/SBOX[8].sbox/t[15] ), .Z(n2424) );
  XOR \b/SBOX[8].sbox/U67  ( .A(\b/SBOX[8].sbox/t[8] ), .B(
        \b/SBOX[8].sbox/t[10] ), .Z(n2425) );
  XOR \b/SBOX[8].sbox/U66  ( .A(\b/SBOX[8].sbox/t[30] ), .B(n2426), .Z(
        \b/SBOX[8].sbox/t[37] ) );
  XOR \b/SBOX[8].sbox/U65  ( .A(\b/SBOX[8].sbox/t[32] ), .B(
        \b/SBOX[8].sbox/t[36] ), .Z(n2426) );
  XOR \b/SBOX[8].sbox/U64  ( .A(msg[71]), .B(msg[66]), .Z(n2446) );
  XOR \b/SBOX[8].sbox/U63  ( .A(\b/SBOX[8].sbox/y[5] ), .B(n2446), .Z(
        \b/SBOX[8].sbox/y[3] ) );
  XOR \b/SBOX[8].sbox/U62  ( .A(n2428), .B(n2427), .Z(\b/SBOX[8].sbox/t[23] )
         );
  XOR \b/SBOX[8].sbox/U61  ( .A(n2430), .B(n2429), .Z(n2427) );
  XOR \b/SBOX[8].sbox/U60  ( .A(n2446), .B(n2431), .Z(n2428) );
  XOR \b/SBOX[8].sbox/U59  ( .A(msg[69]), .B(msg[67]), .Z(n2429) );
  XOR \b/SBOX[8].sbox/U58  ( .A(\b/SBOX[8].sbox/t[12] ), .B(
        \b/SBOX[8].sbox/t[13] ), .Z(n2430) );
  XOR \b/SBOX[8].sbox/U57  ( .A(\b/SBOX[8].sbox/t[7] ), .B(
        \b/SBOX[8].sbox/t[8] ), .Z(n2431) );
  XOR \b/SBOX[8].sbox/U56  ( .A(\b/SBOX[8].sbox/t[36] ), .B(
        \b/SBOX[8].sbox/t[23] ), .Z(\b/SBOX[8].sbox/t[44] ) );
  XOR \b/SBOX[8].sbox/U55  ( .A(n2446), .B(n2432), .Z(\b/SBOX[8].sbox/y[12] )
         );
  XOR \b/SBOX[8].sbox/U54  ( .A(msg[68]), .B(msg[65]), .Z(n2432) );
  XOR \b/SBOX[8].sbox/U53  ( .A(\b/SBOX[8].sbox/y[15] ), .B(n2433), .Z(
        \b/SBOX[8].sbox/y[10] ) );
  XOR \b/SBOX[8].sbox/U52  ( .A(msg[70]), .B(msg[69]), .Z(n2433) );
  XOR \b/SBOX[8].sbox/U51  ( .A(n2446), .B(n2434), .Z(\b/SBOX[8].sbox/y[17] )
         );
  XOR \b/SBOX[8].sbox/U50  ( .A(msg[69]), .B(msg[68]), .Z(n2434) );
  XOR \b/SBOX[8].sbox/U49  ( .A(msg[70]), .B(n2447), .Z(\b/SBOX[8].sbox/y[11] ) );
  XOR \b/SBOX[8].sbox/U48  ( .A(msg[64]), .B(\b/SBOX[8].sbox/y[11] ), .Z(
        \b/SBOX[8].sbox/y[7] ) );
  XOR \b/SBOX[8].sbox/U47  ( .A(msg[64]), .B(\b/SBOX[8].sbox/y[15] ), .Z(
        \b/SBOX[8].sbox/y[6] ) );
  XOR \b/SBOX[8].sbox/U46  ( .A(\b/SBOX[8].sbox/t[26] ), .B(
        \b/SBOX[8].sbox/t[24] ), .Z(\b/SBOX[8].sbox/t[27] ) );
  XOR \b/SBOX[8].sbox/U45  ( .A(\b/SBOX[8].sbox/t[36] ), .B(
        \b/SBOX[8].sbox/t[27] ), .Z(\b/SBOX[8].sbox/t[38] ) );
  XOR \b/SBOX[8].sbox/U44  ( .A(n2448), .B(n2435), .Z(\b/SBOX[8].sbox/t[31] )
         );
  XOR \b/SBOX[8].sbox/U43  ( .A(\b/SBOX[8].sbox/t[26] ), .B(n2449), .Z(n2435)
         );
  XOR \b/SBOX[7].sbox/U157  ( .A(\b/SBOX[7].sbox/z[12] ), .B(n2292), .Z(n2356)
         );
  XOR \b/SBOX[7].sbox/U156  ( .A(\b/SBOX[7].sbox/z[0] ), .B(
        \b/SBOX[7].sbox/z[2] ), .Z(n2292) );
  XOR \b/SBOX[7].sbox/U155  ( .A(n2294), .B(n2293), .Z(n2355) );
  XOR \b/SBOX[7].sbox/U154  ( .A(\b/SBOX[7].sbox/z[15] ), .B(
        \b/SBOX[7].sbox/z[16] ), .Z(n2293) );
  XOR \b/SBOX[7].sbox/U153  ( .A(\b/SBOX[7].sbox/z[5] ), .B(
        \b/SBOX[7].sbox/z[13] ), .Z(n2294) );
  XOR \b/SBOX[7].sbox/U152  ( .A(n2355), .B(n2295), .Z(n2369) );
  XOR \b/SBOX[7].sbox/U151  ( .A(\b/SBOX[7].sbox/z[3] ), .B(n2356), .Z(n2295)
         );
  XOR \b/SBOX[7].sbox/U150  ( .A(n2297), .B(n2296), .Z(n2370) );
  XOR \b/SBOX[7].sbox/U149  ( .A(n2355), .B(n2298), .Z(n2296) );
  XOR \b/SBOX[7].sbox/U148  ( .A(\b/SBOX[7].sbox/z[8] ), .B(
        \b/SBOX[7].sbox/z[12] ), .Z(n2297) );
  XOR \b/SBOX[7].sbox/U147  ( .A(\b/SBOX[7].sbox/z[4] ), .B(
        \b/SBOX[7].sbox/z[7] ), .Z(n2298) );
  XOR \b/SBOX[7].sbox/U146  ( .A(n2356), .B(n2299), .Z(n2358) );
  XOR \b/SBOX[7].sbox/U145  ( .A(\b/SBOX[7].sbox/z[8] ), .B(
        \b/SBOX[7].sbox/z[14] ), .Z(n2299) );
  XOR \b/SBOX[7].sbox/U144  ( .A(n2301), .B(n2300), .Z(n2371) );
  XOR \b/SBOX[7].sbox/U143  ( .A(\b/SBOX[7].sbox/z[17] ), .B(n2358), .Z(n2300)
         );
  XOR \b/SBOX[7].sbox/U142  ( .A(\b/SBOX[7].sbox/z[6] ), .B(
        \b/SBOX[7].sbox/z[15] ), .Z(n2301) );
  XOR \b/SBOX[7].sbox/U141  ( .A(\b/SBOX[7].sbox/z[9] ), .B(n2302), .Z(n2359)
         );
  XOR \b/SBOX[7].sbox/U140  ( .A(\b/SBOX[7].sbox/z[0] ), .B(
        \b/SBOX[7].sbox/z[1] ), .Z(n2302) );
  XOR \b/SBOX[7].sbox/U139  ( .A(\b/SBOX[7].sbox/z[16] ), .B(n2303), .Z(n2357)
         );
  XOR \b/SBOX[7].sbox/U138  ( .A(\b/SBOX[7].sbox/z[10] ), .B(
        \b/SBOX[7].sbox/z[15] ), .Z(n2303) );
  XOR \b/SBOX[7].sbox/U137  ( .A(n2305), .B(n2304), .Z(n2372) );
  XOR \b/SBOX[7].sbox/U136  ( .A(n2359), .B(n2357), .Z(n2304) );
  XOR \b/SBOX[7].sbox/U135  ( .A(\b/SBOX[7].sbox/z[6] ), .B(
        \b/SBOX[7].sbox/z[7] ), .Z(n2305) );
  XOR \b/SBOX[7].sbox/U134  ( .A(\b/SBOX[7].sbox/z[4] ), .B(n2357), .Z(n2360)
         );
  XOR \b/SBOX[7].sbox/U133  ( .A(n2360), .B(n2306), .Z(n2361) );
  XOR \b/SBOX[7].sbox/U132  ( .A(\b/SBOX[7].sbox/z[3] ), .B(
        \b/SBOX[7].sbox/z[7] ), .Z(n2306) );
  XOR \b/SBOX[7].sbox/U131  ( .A(n2358), .B(n2307), .Z(shift_row_out[90]) );
  XOR \b/SBOX[7].sbox/U130  ( .A(\b/SBOX[7].sbox/z[11] ), .B(n2361), .Z(n2307)
         );
  XOR \b/SBOX[7].sbox/U129  ( .A(n2309), .B(n2308), .Z(shift_row_out[91]) );
  XOR \b/SBOX[7].sbox/U128  ( .A(n2360), .B(n2310), .Z(n2308) );
  XOR \b/SBOX[7].sbox/U127  ( .A(\b/SBOX[7].sbox/z[5] ), .B(
        \b/SBOX[7].sbox/z[9] ), .Z(n2309) );
  XOR \b/SBOX[7].sbox/U126  ( .A(\b/SBOX[7].sbox/z[1] ), .B(
        \b/SBOX[7].sbox/z[2] ), .Z(n2310) );
  XOR \b/SBOX[7].sbox/U125  ( .A(n2359), .B(n2311), .Z(shift_row_out[92]) );
  XOR \b/SBOX[7].sbox/U124  ( .A(\b/SBOX[7].sbox/z[3] ), .B(n2360), .Z(n2311)
         );
  XOR \b/SBOX[7].sbox/U123  ( .A(n2361), .B(n2312), .Z(shift_row_out[95]) );
  XOR \b/SBOX[7].sbox/U122  ( .A(\b/SBOX[7].sbox/z[6] ), .B(
        \b/SBOX[7].sbox/z[9] ), .Z(n2312) );
  XOR \b/SBOX[7].sbox/U121  ( .A(n2314), .B(n2313), .Z(n2362) );
  XOR \b/SBOX[7].sbox/U120  ( .A(n2316), .B(n2315), .Z(n2313) );
  XOR \b/SBOX[7].sbox/U119  ( .A(msg[61]), .B(msg[57]), .Z(n2314) );
  XOR \b/SBOX[7].sbox/U118  ( .A(\b/SBOX[7].sbox/t[36] ), .B(
        \b/SBOX[7].sbox/t[39] ), .Z(n2315) );
  XOR \b/SBOX[7].sbox/U117  ( .A(\b/SBOX[7].sbox/t[3] ), .B(
        \b/SBOX[7].sbox/t[8] ), .Z(n2316) );
  XOR \b/SBOX[7].sbox/U116  ( .A(n2318), .B(n2317), .Z(\b/SBOX[7].sbox/t[41] )
         );
  XOR \b/SBOX[7].sbox/U115  ( .A(n2362), .B(n2319), .Z(n2317) );
  XOR \b/SBOX[7].sbox/U114  ( .A(\b/SBOX[7].sbox/t[32] ), .B(msg[63]), .Z(
        n2318) );
  XOR \b/SBOX[7].sbox/U113  ( .A(\b/SBOX[7].sbox/t[5] ), .B(
        \b/SBOX[7].sbox/t[10] ), .Z(n2319) );
  XOR \b/SBOX[7].sbox/U112  ( .A(\b/SBOX[7].sbox/t[2] ), .B(msg[62]), .Z(n2363) );
  XOR \b/SBOX[7].sbox/U111  ( .A(n2321), .B(n2320), .Z(\b/SBOX[7].sbox/t[45] )
         );
  XOR \b/SBOX[7].sbox/U110  ( .A(n2363), .B(n2322), .Z(n2320) );
  XOR \b/SBOX[7].sbox/U109  ( .A(msg[60]), .B(n2362), .Z(n2321) );
  XOR \b/SBOX[7].sbox/U108  ( .A(\b/SBOX[7].sbox/t[7] ), .B(
        \b/SBOX[7].sbox/t[28] ), .Z(n2322) );
  XOR \b/SBOX[7].sbox/U107  ( .A(n2363), .B(n2323), .Z(n2368) );
  XOR \b/SBOX[7].sbox/U106  ( .A(\b/SBOX[7].sbox/t[5] ), .B(msg[60]), .Z(n2323) );
  XOR \b/SBOX[7].sbox/U105  ( .A(msg[63]), .B(n2324), .Z(n2364) );
  XOR \b/SBOX[7].sbox/U104  ( .A(\b/SBOX[7].sbox/t[7] ), .B(
        \b/SBOX[7].sbox/t[10] ), .Z(n2324) );
  XOR \b/SBOX[7].sbox/U103  ( .A(n2326), .B(n2325), .Z(\b/SBOX[7].sbox/t[42] )
         );
  XOR \b/SBOX[7].sbox/U102  ( .A(n2368), .B(n2364), .Z(n2325) );
  XOR \b/SBOX[7].sbox/U101  ( .A(\b/SBOX[7].sbox/t[28] ), .B(
        \b/SBOX[7].sbox/t[32] ), .Z(n2326) );
  XOR \b/SBOX[7].sbox/U100  ( .A(msg[57]), .B(n2327), .Z(n2366) );
  XOR \b/SBOX[7].sbox/U99  ( .A(msg[59]), .B(msg[58]), .Z(n2327) );
  XOR \b/SBOX[7].sbox/U98  ( .A(msg[61]), .B(n2366), .Z(\b/SBOX[7].sbox/y[16] ) );
  XOR \b/SBOX[7].sbox/U97  ( .A(\b/SBOX[7].sbox/y[16] ), .B(n2328), .Z(n2367)
         );
  XOR \b/SBOX[7].sbox/U96  ( .A(\b/SBOX[7].sbox/t[12] ), .B(
        \b/SBOX[7].sbox/t[15] ), .Z(n2328) );
  XOR \b/SBOX[7].sbox/U95  ( .A(n2367), .B(n2329), .Z(\b/SBOX[7].sbox/t[29] )
         );
  XOR \b/SBOX[7].sbox/U94  ( .A(\b/SBOX[7].sbox/t[28] ), .B(n2368), .Z(n2329)
         );
  XOR \b/SBOX[7].sbox/U93  ( .A(msg[56]), .B(n2330), .Z(\b/SBOX[7].sbox/y[1] )
         );
  XOR \b/SBOX[7].sbox/U92  ( .A(msg[62]), .B(msg[61]), .Z(n2330) );
  XOR \b/SBOX[7].sbox/U91  ( .A(msg[63]), .B(\b/SBOX[7].sbox/y[1] ), .Z(
        \b/SBOX[7].sbox/y[2] ) );
  XOR \b/SBOX[7].sbox/U90  ( .A(n2332), .B(n2331), .Z(\b/SBOX[7].sbox/t[25] )
         );
  XOR \b/SBOX[7].sbox/U89  ( .A(n2334), .B(n2333), .Z(n2331) );
  XOR \b/SBOX[7].sbox/U88  ( .A(msg[63]), .B(msg[61]), .Z(n2332) );
  XOR \b/SBOX[7].sbox/U87  ( .A(\b/SBOX[7].sbox/t[13] ), .B(
        \b/SBOX[7].sbox/t[15] ), .Z(n2333) );
  XOR \b/SBOX[7].sbox/U86  ( .A(\b/SBOX[7].sbox/t[3] ), .B(
        \b/SBOX[7].sbox/t[5] ), .Z(n2334) );
  XOR \b/SBOX[7].sbox/U85  ( .A(\b/SBOX[7].sbox/t[39] ), .B(
        \b/SBOX[7].sbox/t[25] ), .Z(\b/SBOX[7].sbox/t[40] ) );
  XOR \b/SBOX[7].sbox/U84  ( .A(msg[57]), .B(\b/SBOX[7].sbox/y[1] ), .Z(
        \b/SBOX[7].sbox/y[5] ) );
  XOR \b/SBOX[7].sbox/U83  ( .A(n2336), .B(n2335), .Z(\b/SBOX[7].sbox/y[15] )
         );
  XOR \b/SBOX[7].sbox/U82  ( .A(msg[59]), .B(msg[57]), .Z(n2335) );
  XOR \b/SBOX[7].sbox/U81  ( .A(msg[63]), .B(msg[60]), .Z(n2336) );
  XOR \b/SBOX[7].sbox/U80  ( .A(n2338), .B(n2337), .Z(\b/SBOX[7].sbox/t[21] )
         );
  XOR \b/SBOX[7].sbox/U79  ( .A(n2340), .B(n2339), .Z(n2337) );
  XOR \b/SBOX[7].sbox/U78  ( .A(\b/SBOX[7].sbox/y[15] ), .B(n2363), .Z(n2338)
         );
  XOR \b/SBOX[7].sbox/U77  ( .A(\b/SBOX[7].sbox/t[13] ), .B(msg[58]), .Z(n2339) );
  XOR \b/SBOX[7].sbox/U76  ( .A(\b/SBOX[7].sbox/t[3] ), .B(
        \b/SBOX[7].sbox/t[12] ), .Z(n2340) );
  XOR \b/SBOX[7].sbox/U75  ( .A(\b/SBOX[7].sbox/t[21] ), .B(n2341), .Z(
        \b/SBOX[7].sbox/t[43] ) );
  XOR \b/SBOX[7].sbox/U74  ( .A(\b/SBOX[7].sbox/t[28] ), .B(
        \b/SBOX[7].sbox/t[39] ), .Z(n2341) );
  XOR \b/SBOX[7].sbox/U73  ( .A(n2367), .B(n2364), .Z(\b/SBOX[7].sbox/t[24] )
         );
  XOR \b/SBOX[7].sbox/U72  ( .A(\b/SBOX[7].sbox/t[32] ), .B(
        \b/SBOX[7].sbox/t[24] ), .Z(\b/SBOX[7].sbox/t[33] ) );
  XOR \b/SBOX[7].sbox/U71  ( .A(msg[60]), .B(\b/SBOX[7].sbox/y[1] ), .Z(
        \b/SBOX[7].sbox/y[4] ) );
  XOR \b/SBOX[7].sbox/U70  ( .A(n2343), .B(n2342), .Z(\b/SBOX[7].sbox/t[30] )
         );
  XOR \b/SBOX[7].sbox/U69  ( .A(msg[57]), .B(n2344), .Z(n2342) );
  XOR \b/SBOX[7].sbox/U68  ( .A(\b/SBOX[7].sbox/t[13] ), .B(
        \b/SBOX[7].sbox/t[15] ), .Z(n2343) );
  XOR \b/SBOX[7].sbox/U67  ( .A(\b/SBOX[7].sbox/t[8] ), .B(
        \b/SBOX[7].sbox/t[10] ), .Z(n2344) );
  XOR \b/SBOX[7].sbox/U66  ( .A(\b/SBOX[7].sbox/t[30] ), .B(n2345), .Z(
        \b/SBOX[7].sbox/t[37] ) );
  XOR \b/SBOX[7].sbox/U65  ( .A(\b/SBOX[7].sbox/t[32] ), .B(
        \b/SBOX[7].sbox/t[36] ), .Z(n2345) );
  XOR \b/SBOX[7].sbox/U64  ( .A(msg[63]), .B(msg[58]), .Z(n2365) );
  XOR \b/SBOX[7].sbox/U63  ( .A(\b/SBOX[7].sbox/y[5] ), .B(n2365), .Z(
        \b/SBOX[7].sbox/y[3] ) );
  XOR \b/SBOX[7].sbox/U62  ( .A(n2347), .B(n2346), .Z(\b/SBOX[7].sbox/t[23] )
         );
  XOR \b/SBOX[7].sbox/U61  ( .A(n2349), .B(n2348), .Z(n2346) );
  XOR \b/SBOX[7].sbox/U60  ( .A(n2365), .B(n2350), .Z(n2347) );
  XOR \b/SBOX[7].sbox/U59  ( .A(msg[61]), .B(msg[59]), .Z(n2348) );
  XOR \b/SBOX[7].sbox/U58  ( .A(\b/SBOX[7].sbox/t[12] ), .B(
        \b/SBOX[7].sbox/t[13] ), .Z(n2349) );
  XOR \b/SBOX[7].sbox/U57  ( .A(\b/SBOX[7].sbox/t[7] ), .B(
        \b/SBOX[7].sbox/t[8] ), .Z(n2350) );
  XOR \b/SBOX[7].sbox/U56  ( .A(\b/SBOX[7].sbox/t[36] ), .B(
        \b/SBOX[7].sbox/t[23] ), .Z(\b/SBOX[7].sbox/t[44] ) );
  XOR \b/SBOX[7].sbox/U55  ( .A(n2365), .B(n2351), .Z(\b/SBOX[7].sbox/y[12] )
         );
  XOR \b/SBOX[7].sbox/U54  ( .A(msg[60]), .B(msg[57]), .Z(n2351) );
  XOR \b/SBOX[7].sbox/U53  ( .A(\b/SBOX[7].sbox/y[15] ), .B(n2352), .Z(
        \b/SBOX[7].sbox/y[10] ) );
  XOR \b/SBOX[7].sbox/U52  ( .A(msg[62]), .B(msg[61]), .Z(n2352) );
  XOR \b/SBOX[7].sbox/U51  ( .A(n2365), .B(n2353), .Z(\b/SBOX[7].sbox/y[17] )
         );
  XOR \b/SBOX[7].sbox/U50  ( .A(msg[61]), .B(msg[60]), .Z(n2353) );
  XOR \b/SBOX[7].sbox/U49  ( .A(msg[62]), .B(n2366), .Z(\b/SBOX[7].sbox/y[11] ) );
  XOR \b/SBOX[7].sbox/U48  ( .A(msg[56]), .B(\b/SBOX[7].sbox/y[11] ), .Z(
        \b/SBOX[7].sbox/y[7] ) );
  XOR \b/SBOX[7].sbox/U47  ( .A(msg[56]), .B(\b/SBOX[7].sbox/y[15] ), .Z(
        \b/SBOX[7].sbox/y[6] ) );
  XOR \b/SBOX[7].sbox/U46  ( .A(\b/SBOX[7].sbox/t[26] ), .B(
        \b/SBOX[7].sbox/t[24] ), .Z(\b/SBOX[7].sbox/t[27] ) );
  XOR \b/SBOX[7].sbox/U45  ( .A(\b/SBOX[7].sbox/t[36] ), .B(
        \b/SBOX[7].sbox/t[27] ), .Z(\b/SBOX[7].sbox/t[38] ) );
  XOR \b/SBOX[7].sbox/U44  ( .A(n2367), .B(n2354), .Z(\b/SBOX[7].sbox/t[31] )
         );
  XOR \b/SBOX[7].sbox/U43  ( .A(\b/SBOX[7].sbox/t[26] ), .B(n2368), .Z(n2354)
         );
  XOR \b/SBOX[6].sbox/U157  ( .A(\b/SBOX[6].sbox/z[12] ), .B(n2211), .Z(n2275)
         );
  XOR \b/SBOX[6].sbox/U156  ( .A(\b/SBOX[6].sbox/z[0] ), .B(
        \b/SBOX[6].sbox/z[2] ), .Z(n2211) );
  XOR \b/SBOX[6].sbox/U155  ( .A(n2213), .B(n2212), .Z(n2274) );
  XOR \b/SBOX[6].sbox/U154  ( .A(\b/SBOX[6].sbox/z[15] ), .B(
        \b/SBOX[6].sbox/z[16] ), .Z(n2212) );
  XOR \b/SBOX[6].sbox/U153  ( .A(\b/SBOX[6].sbox/z[5] ), .B(
        \b/SBOX[6].sbox/z[13] ), .Z(n2213) );
  XOR \b/SBOX[6].sbox/U152  ( .A(n2274), .B(n2214), .Z(n2288) );
  XOR \b/SBOX[6].sbox/U151  ( .A(\b/SBOX[6].sbox/z[3] ), .B(n2275), .Z(n2214)
         );
  XOR \b/SBOX[6].sbox/U150  ( .A(n2216), .B(n2215), .Z(n2289) );
  XOR \b/SBOX[6].sbox/U149  ( .A(n2274), .B(n2217), .Z(n2215) );
  XOR \b/SBOX[6].sbox/U148  ( .A(\b/SBOX[6].sbox/z[8] ), .B(
        \b/SBOX[6].sbox/z[12] ), .Z(n2216) );
  XOR \b/SBOX[6].sbox/U147  ( .A(\b/SBOX[6].sbox/z[4] ), .B(
        \b/SBOX[6].sbox/z[7] ), .Z(n2217) );
  XOR \b/SBOX[6].sbox/U146  ( .A(n2275), .B(n2218), .Z(n2277) );
  XOR \b/SBOX[6].sbox/U145  ( .A(\b/SBOX[6].sbox/z[8] ), .B(
        \b/SBOX[6].sbox/z[14] ), .Z(n2218) );
  XOR \b/SBOX[6].sbox/U144  ( .A(n2220), .B(n2219), .Z(n2290) );
  XOR \b/SBOX[6].sbox/U143  ( .A(\b/SBOX[6].sbox/z[17] ), .B(n2277), .Z(n2219)
         );
  XOR \b/SBOX[6].sbox/U142  ( .A(\b/SBOX[6].sbox/z[6] ), .B(
        \b/SBOX[6].sbox/z[15] ), .Z(n2220) );
  XOR \b/SBOX[6].sbox/U141  ( .A(\b/SBOX[6].sbox/z[9] ), .B(n2221), .Z(n2278)
         );
  XOR \b/SBOX[6].sbox/U140  ( .A(\b/SBOX[6].sbox/z[0] ), .B(
        \b/SBOX[6].sbox/z[1] ), .Z(n2221) );
  XOR \b/SBOX[6].sbox/U139  ( .A(\b/SBOX[6].sbox/z[16] ), .B(n2222), .Z(n2276)
         );
  XOR \b/SBOX[6].sbox/U138  ( .A(\b/SBOX[6].sbox/z[10] ), .B(
        \b/SBOX[6].sbox/z[15] ), .Z(n2222) );
  XOR \b/SBOX[6].sbox/U137  ( .A(n2224), .B(n2223), .Z(n2291) );
  XOR \b/SBOX[6].sbox/U136  ( .A(n2278), .B(n2276), .Z(n2223) );
  XOR \b/SBOX[6].sbox/U135  ( .A(\b/SBOX[6].sbox/z[6] ), .B(
        \b/SBOX[6].sbox/z[7] ), .Z(n2224) );
  XOR \b/SBOX[6].sbox/U134  ( .A(\b/SBOX[6].sbox/z[4] ), .B(n2276), .Z(n2279)
         );
  XOR \b/SBOX[6].sbox/U133  ( .A(n2279), .B(n2225), .Z(n2280) );
  XOR \b/SBOX[6].sbox/U132  ( .A(\b/SBOX[6].sbox/z[3] ), .B(
        \b/SBOX[6].sbox/z[7] ), .Z(n2225) );
  XOR \b/SBOX[6].sbox/U131  ( .A(n2277), .B(n2226), .Z(shift_row_out[114]) );
  XOR \b/SBOX[6].sbox/U130  ( .A(\b/SBOX[6].sbox/z[11] ), .B(n2280), .Z(n2226)
         );
  XOR \b/SBOX[6].sbox/U129  ( .A(n2228), .B(n2227), .Z(shift_row_out[115]) );
  XOR \b/SBOX[6].sbox/U128  ( .A(n2279), .B(n2229), .Z(n2227) );
  XOR \b/SBOX[6].sbox/U127  ( .A(\b/SBOX[6].sbox/z[5] ), .B(
        \b/SBOX[6].sbox/z[9] ), .Z(n2228) );
  XOR \b/SBOX[6].sbox/U126  ( .A(\b/SBOX[6].sbox/z[1] ), .B(
        \b/SBOX[6].sbox/z[2] ), .Z(n2229) );
  XOR \b/SBOX[6].sbox/U125  ( .A(n2278), .B(n2230), .Z(shift_row_out[116]) );
  XOR \b/SBOX[6].sbox/U124  ( .A(\b/SBOX[6].sbox/z[3] ), .B(n2279), .Z(n2230)
         );
  XOR \b/SBOX[6].sbox/U123  ( .A(n2280), .B(n2231), .Z(shift_row_out[119]) );
  XOR \b/SBOX[6].sbox/U122  ( .A(\b/SBOX[6].sbox/z[6] ), .B(
        \b/SBOX[6].sbox/z[9] ), .Z(n2231) );
  XOR \b/SBOX[6].sbox/U121  ( .A(n2233), .B(n2232), .Z(n2281) );
  XOR \b/SBOX[6].sbox/U120  ( .A(n2235), .B(n2234), .Z(n2232) );
  XOR \b/SBOX[6].sbox/U119  ( .A(msg[53]), .B(msg[49]), .Z(n2233) );
  XOR \b/SBOX[6].sbox/U118  ( .A(\b/SBOX[6].sbox/t[36] ), .B(
        \b/SBOX[6].sbox/t[39] ), .Z(n2234) );
  XOR \b/SBOX[6].sbox/U117  ( .A(\b/SBOX[6].sbox/t[3] ), .B(
        \b/SBOX[6].sbox/t[8] ), .Z(n2235) );
  XOR \b/SBOX[6].sbox/U116  ( .A(n2237), .B(n2236), .Z(\b/SBOX[6].sbox/t[41] )
         );
  XOR \b/SBOX[6].sbox/U115  ( .A(n2281), .B(n2238), .Z(n2236) );
  XOR \b/SBOX[6].sbox/U114  ( .A(\b/SBOX[6].sbox/t[32] ), .B(msg[55]), .Z(
        n2237) );
  XOR \b/SBOX[6].sbox/U113  ( .A(\b/SBOX[6].sbox/t[5] ), .B(
        \b/SBOX[6].sbox/t[10] ), .Z(n2238) );
  XOR \b/SBOX[6].sbox/U112  ( .A(\b/SBOX[6].sbox/t[2] ), .B(msg[54]), .Z(n2282) );
  XOR \b/SBOX[6].sbox/U111  ( .A(n2240), .B(n2239), .Z(\b/SBOX[6].sbox/t[45] )
         );
  XOR \b/SBOX[6].sbox/U110  ( .A(n2282), .B(n2241), .Z(n2239) );
  XOR \b/SBOX[6].sbox/U109  ( .A(msg[52]), .B(n2281), .Z(n2240) );
  XOR \b/SBOX[6].sbox/U108  ( .A(\b/SBOX[6].sbox/t[7] ), .B(
        \b/SBOX[6].sbox/t[28] ), .Z(n2241) );
  XOR \b/SBOX[6].sbox/U107  ( .A(n2282), .B(n2242), .Z(n2287) );
  XOR \b/SBOX[6].sbox/U106  ( .A(\b/SBOX[6].sbox/t[5] ), .B(msg[52]), .Z(n2242) );
  XOR \b/SBOX[6].sbox/U105  ( .A(msg[55]), .B(n2243), .Z(n2283) );
  XOR \b/SBOX[6].sbox/U104  ( .A(\b/SBOX[6].sbox/t[7] ), .B(
        \b/SBOX[6].sbox/t[10] ), .Z(n2243) );
  XOR \b/SBOX[6].sbox/U103  ( .A(n2245), .B(n2244), .Z(\b/SBOX[6].sbox/t[42] )
         );
  XOR \b/SBOX[6].sbox/U102  ( .A(n2287), .B(n2283), .Z(n2244) );
  XOR \b/SBOX[6].sbox/U101  ( .A(\b/SBOX[6].sbox/t[28] ), .B(
        \b/SBOX[6].sbox/t[32] ), .Z(n2245) );
  XOR \b/SBOX[6].sbox/U100  ( .A(msg[49]), .B(n2246), .Z(n2285) );
  XOR \b/SBOX[6].sbox/U99  ( .A(msg[51]), .B(msg[50]), .Z(n2246) );
  XOR \b/SBOX[6].sbox/U98  ( .A(msg[53]), .B(n2285), .Z(\b/SBOX[6].sbox/y[16] ) );
  XOR \b/SBOX[6].sbox/U97  ( .A(\b/SBOX[6].sbox/y[16] ), .B(n2247), .Z(n2286)
         );
  XOR \b/SBOX[6].sbox/U96  ( .A(\b/SBOX[6].sbox/t[12] ), .B(
        \b/SBOX[6].sbox/t[15] ), .Z(n2247) );
  XOR \b/SBOX[6].sbox/U95  ( .A(n2286), .B(n2248), .Z(\b/SBOX[6].sbox/t[29] )
         );
  XOR \b/SBOX[6].sbox/U94  ( .A(\b/SBOX[6].sbox/t[28] ), .B(n2287), .Z(n2248)
         );
  XOR \b/SBOX[6].sbox/U93  ( .A(msg[48]), .B(n2249), .Z(\b/SBOX[6].sbox/y[1] )
         );
  XOR \b/SBOX[6].sbox/U92  ( .A(msg[54]), .B(msg[53]), .Z(n2249) );
  XOR \b/SBOX[6].sbox/U91  ( .A(msg[55]), .B(\b/SBOX[6].sbox/y[1] ), .Z(
        \b/SBOX[6].sbox/y[2] ) );
  XOR \b/SBOX[6].sbox/U90  ( .A(n2251), .B(n2250), .Z(\b/SBOX[6].sbox/t[25] )
         );
  XOR \b/SBOX[6].sbox/U89  ( .A(n2253), .B(n2252), .Z(n2250) );
  XOR \b/SBOX[6].sbox/U88  ( .A(msg[55]), .B(msg[53]), .Z(n2251) );
  XOR \b/SBOX[6].sbox/U87  ( .A(\b/SBOX[6].sbox/t[13] ), .B(
        \b/SBOX[6].sbox/t[15] ), .Z(n2252) );
  XOR \b/SBOX[6].sbox/U86  ( .A(\b/SBOX[6].sbox/t[3] ), .B(
        \b/SBOX[6].sbox/t[5] ), .Z(n2253) );
  XOR \b/SBOX[6].sbox/U85  ( .A(\b/SBOX[6].sbox/t[39] ), .B(
        \b/SBOX[6].sbox/t[25] ), .Z(\b/SBOX[6].sbox/t[40] ) );
  XOR \b/SBOX[6].sbox/U84  ( .A(msg[49]), .B(\b/SBOX[6].sbox/y[1] ), .Z(
        \b/SBOX[6].sbox/y[5] ) );
  XOR \b/SBOX[6].sbox/U83  ( .A(n2255), .B(n2254), .Z(\b/SBOX[6].sbox/y[15] )
         );
  XOR \b/SBOX[6].sbox/U82  ( .A(msg[51]), .B(msg[49]), .Z(n2254) );
  XOR \b/SBOX[6].sbox/U81  ( .A(msg[55]), .B(msg[52]), .Z(n2255) );
  XOR \b/SBOX[6].sbox/U80  ( .A(n2257), .B(n2256), .Z(\b/SBOX[6].sbox/t[21] )
         );
  XOR \b/SBOX[6].sbox/U79  ( .A(n2259), .B(n2258), .Z(n2256) );
  XOR \b/SBOX[6].sbox/U78  ( .A(\b/SBOX[6].sbox/y[15] ), .B(n2282), .Z(n2257)
         );
  XOR \b/SBOX[6].sbox/U77  ( .A(\b/SBOX[6].sbox/t[13] ), .B(msg[50]), .Z(n2258) );
  XOR \b/SBOX[6].sbox/U76  ( .A(\b/SBOX[6].sbox/t[3] ), .B(
        \b/SBOX[6].sbox/t[12] ), .Z(n2259) );
  XOR \b/SBOX[6].sbox/U75  ( .A(\b/SBOX[6].sbox/t[21] ), .B(n2260), .Z(
        \b/SBOX[6].sbox/t[43] ) );
  XOR \b/SBOX[6].sbox/U74  ( .A(\b/SBOX[6].sbox/t[28] ), .B(
        \b/SBOX[6].sbox/t[39] ), .Z(n2260) );
  XOR \b/SBOX[6].sbox/U73  ( .A(n2286), .B(n2283), .Z(\b/SBOX[6].sbox/t[24] )
         );
  XOR \b/SBOX[6].sbox/U72  ( .A(\b/SBOX[6].sbox/t[32] ), .B(
        \b/SBOX[6].sbox/t[24] ), .Z(\b/SBOX[6].sbox/t[33] ) );
  XOR \b/SBOX[6].sbox/U71  ( .A(msg[52]), .B(\b/SBOX[6].sbox/y[1] ), .Z(
        \b/SBOX[6].sbox/y[4] ) );
  XOR \b/SBOX[6].sbox/U70  ( .A(n2262), .B(n2261), .Z(\b/SBOX[6].sbox/t[30] )
         );
  XOR \b/SBOX[6].sbox/U69  ( .A(msg[49]), .B(n2263), .Z(n2261) );
  XOR \b/SBOX[6].sbox/U68  ( .A(\b/SBOX[6].sbox/t[13] ), .B(
        \b/SBOX[6].sbox/t[15] ), .Z(n2262) );
  XOR \b/SBOX[6].sbox/U67  ( .A(\b/SBOX[6].sbox/t[8] ), .B(
        \b/SBOX[6].sbox/t[10] ), .Z(n2263) );
  XOR \b/SBOX[6].sbox/U66  ( .A(\b/SBOX[6].sbox/t[30] ), .B(n2264), .Z(
        \b/SBOX[6].sbox/t[37] ) );
  XOR \b/SBOX[6].sbox/U65  ( .A(\b/SBOX[6].sbox/t[32] ), .B(
        \b/SBOX[6].sbox/t[36] ), .Z(n2264) );
  XOR \b/SBOX[6].sbox/U64  ( .A(msg[55]), .B(msg[50]), .Z(n2284) );
  XOR \b/SBOX[6].sbox/U63  ( .A(\b/SBOX[6].sbox/y[5] ), .B(n2284), .Z(
        \b/SBOX[6].sbox/y[3] ) );
  XOR \b/SBOX[6].sbox/U62  ( .A(n2266), .B(n2265), .Z(\b/SBOX[6].sbox/t[23] )
         );
  XOR \b/SBOX[6].sbox/U61  ( .A(n2268), .B(n2267), .Z(n2265) );
  XOR \b/SBOX[6].sbox/U60  ( .A(n2284), .B(n2269), .Z(n2266) );
  XOR \b/SBOX[6].sbox/U59  ( .A(msg[53]), .B(msg[51]), .Z(n2267) );
  XOR \b/SBOX[6].sbox/U58  ( .A(\b/SBOX[6].sbox/t[12] ), .B(
        \b/SBOX[6].sbox/t[13] ), .Z(n2268) );
  XOR \b/SBOX[6].sbox/U57  ( .A(\b/SBOX[6].sbox/t[7] ), .B(
        \b/SBOX[6].sbox/t[8] ), .Z(n2269) );
  XOR \b/SBOX[6].sbox/U56  ( .A(\b/SBOX[6].sbox/t[36] ), .B(
        \b/SBOX[6].sbox/t[23] ), .Z(\b/SBOX[6].sbox/t[44] ) );
  XOR \b/SBOX[6].sbox/U55  ( .A(n2284), .B(n2270), .Z(\b/SBOX[6].sbox/y[12] )
         );
  XOR \b/SBOX[6].sbox/U54  ( .A(msg[52]), .B(msg[49]), .Z(n2270) );
  XOR \b/SBOX[6].sbox/U53  ( .A(\b/SBOX[6].sbox/y[15] ), .B(n2271), .Z(
        \b/SBOX[6].sbox/y[10] ) );
  XOR \b/SBOX[6].sbox/U52  ( .A(msg[54]), .B(msg[53]), .Z(n2271) );
  XOR \b/SBOX[6].sbox/U51  ( .A(n2284), .B(n2272), .Z(\b/SBOX[6].sbox/y[17] )
         );
  XOR \b/SBOX[6].sbox/U50  ( .A(msg[53]), .B(msg[52]), .Z(n2272) );
  XOR \b/SBOX[6].sbox/U49  ( .A(msg[54]), .B(n2285), .Z(\b/SBOX[6].sbox/y[11] ) );
  XOR \b/SBOX[6].sbox/U48  ( .A(msg[48]), .B(\b/SBOX[6].sbox/y[11] ), .Z(
        \b/SBOX[6].sbox/y[7] ) );
  XOR \b/SBOX[6].sbox/U47  ( .A(msg[48]), .B(\b/SBOX[6].sbox/y[15] ), .Z(
        \b/SBOX[6].sbox/y[6] ) );
  XOR \b/SBOX[6].sbox/U46  ( .A(\b/SBOX[6].sbox/t[26] ), .B(
        \b/SBOX[6].sbox/t[24] ), .Z(\b/SBOX[6].sbox/t[27] ) );
  XOR \b/SBOX[6].sbox/U45  ( .A(\b/SBOX[6].sbox/t[36] ), .B(
        \b/SBOX[6].sbox/t[27] ), .Z(\b/SBOX[6].sbox/t[38] ) );
  XOR \b/SBOX[6].sbox/U44  ( .A(n2286), .B(n2273), .Z(\b/SBOX[6].sbox/t[31] )
         );
  XOR \b/SBOX[6].sbox/U43  ( .A(\b/SBOX[6].sbox/t[26] ), .B(n2287), .Z(n2273)
         );
  XOR \b/SBOX[5].sbox/U157  ( .A(\b/SBOX[5].sbox/z[12] ), .B(n2130), .Z(n2194)
         );
  XOR \b/SBOX[5].sbox/U156  ( .A(\b/SBOX[5].sbox/z[0] ), .B(
        \b/SBOX[5].sbox/z[2] ), .Z(n2130) );
  XOR \b/SBOX[5].sbox/U155  ( .A(n2132), .B(n2131), .Z(n2193) );
  XOR \b/SBOX[5].sbox/U154  ( .A(\b/SBOX[5].sbox/z[15] ), .B(
        \b/SBOX[5].sbox/z[16] ), .Z(n2131) );
  XOR \b/SBOX[5].sbox/U153  ( .A(\b/SBOX[5].sbox/z[5] ), .B(
        \b/SBOX[5].sbox/z[13] ), .Z(n2132) );
  XOR \b/SBOX[5].sbox/U152  ( .A(n2193), .B(n2133), .Z(n2207) );
  XOR \b/SBOX[5].sbox/U151  ( .A(\b/SBOX[5].sbox/z[3] ), .B(n2194), .Z(n2133)
         );
  XOR \b/SBOX[5].sbox/U150  ( .A(n2135), .B(n2134), .Z(n2208) );
  XOR \b/SBOX[5].sbox/U149  ( .A(n2193), .B(n2136), .Z(n2134) );
  XOR \b/SBOX[5].sbox/U148  ( .A(\b/SBOX[5].sbox/z[8] ), .B(
        \b/SBOX[5].sbox/z[12] ), .Z(n2135) );
  XOR \b/SBOX[5].sbox/U147  ( .A(\b/SBOX[5].sbox/z[4] ), .B(
        \b/SBOX[5].sbox/z[7] ), .Z(n2136) );
  XOR \b/SBOX[5].sbox/U146  ( .A(n2194), .B(n2137), .Z(n2196) );
  XOR \b/SBOX[5].sbox/U145  ( .A(\b/SBOX[5].sbox/z[8] ), .B(
        \b/SBOX[5].sbox/z[14] ), .Z(n2137) );
  XOR \b/SBOX[5].sbox/U144  ( .A(n2139), .B(n2138), .Z(n2209) );
  XOR \b/SBOX[5].sbox/U143  ( .A(\b/SBOX[5].sbox/z[17] ), .B(n2196), .Z(n2138)
         );
  XOR \b/SBOX[5].sbox/U142  ( .A(\b/SBOX[5].sbox/z[6] ), .B(
        \b/SBOX[5].sbox/z[15] ), .Z(n2139) );
  XOR \b/SBOX[5].sbox/U141  ( .A(\b/SBOX[5].sbox/z[9] ), .B(n2140), .Z(n2197)
         );
  XOR \b/SBOX[5].sbox/U140  ( .A(\b/SBOX[5].sbox/z[0] ), .B(
        \b/SBOX[5].sbox/z[1] ), .Z(n2140) );
  XOR \b/SBOX[5].sbox/U139  ( .A(\b/SBOX[5].sbox/z[16] ), .B(n2141), .Z(n2195)
         );
  XOR \b/SBOX[5].sbox/U138  ( .A(\b/SBOX[5].sbox/z[10] ), .B(
        \b/SBOX[5].sbox/z[15] ), .Z(n2141) );
  XOR \b/SBOX[5].sbox/U137  ( .A(n2143), .B(n2142), .Z(n2210) );
  XOR \b/SBOX[5].sbox/U136  ( .A(n2197), .B(n2195), .Z(n2142) );
  XOR \b/SBOX[5].sbox/U135  ( .A(\b/SBOX[5].sbox/z[6] ), .B(
        \b/SBOX[5].sbox/z[7] ), .Z(n2143) );
  XOR \b/SBOX[5].sbox/U134  ( .A(\b/SBOX[5].sbox/z[4] ), .B(n2195), .Z(n2198)
         );
  XOR \b/SBOX[5].sbox/U133  ( .A(n2198), .B(n2144), .Z(n2199) );
  XOR \b/SBOX[5].sbox/U132  ( .A(\b/SBOX[5].sbox/z[3] ), .B(
        \b/SBOX[5].sbox/z[7] ), .Z(n2144) );
  XOR \b/SBOX[5].sbox/U131  ( .A(n2196), .B(n2145), .Z(shift_row_out[10]) );
  XOR \b/SBOX[5].sbox/U130  ( .A(\b/SBOX[5].sbox/z[11] ), .B(n2199), .Z(n2145)
         );
  XOR \b/SBOX[5].sbox/U129  ( .A(n2147), .B(n2146), .Z(shift_row_out[11]) );
  XOR \b/SBOX[5].sbox/U128  ( .A(n2198), .B(n2148), .Z(n2146) );
  XOR \b/SBOX[5].sbox/U127  ( .A(\b/SBOX[5].sbox/z[5] ), .B(
        \b/SBOX[5].sbox/z[9] ), .Z(n2147) );
  XOR \b/SBOX[5].sbox/U126  ( .A(\b/SBOX[5].sbox/z[1] ), .B(
        \b/SBOX[5].sbox/z[2] ), .Z(n2148) );
  XOR \b/SBOX[5].sbox/U125  ( .A(n2197), .B(n2149), .Z(shift_row_out[12]) );
  XOR \b/SBOX[5].sbox/U124  ( .A(\b/SBOX[5].sbox/z[3] ), .B(n2198), .Z(n2149)
         );
  XOR \b/SBOX[5].sbox/U123  ( .A(n2199), .B(n2150), .Z(shift_row_out[15]) );
  XOR \b/SBOX[5].sbox/U122  ( .A(\b/SBOX[5].sbox/z[6] ), .B(
        \b/SBOX[5].sbox/z[9] ), .Z(n2150) );
  XOR \b/SBOX[5].sbox/U121  ( .A(n2152), .B(n2151), .Z(n2200) );
  XOR \b/SBOX[5].sbox/U120  ( .A(n2154), .B(n2153), .Z(n2151) );
  XOR \b/SBOX[5].sbox/U119  ( .A(msg[45]), .B(msg[41]), .Z(n2152) );
  XOR \b/SBOX[5].sbox/U118  ( .A(\b/SBOX[5].sbox/t[36] ), .B(
        \b/SBOX[5].sbox/t[39] ), .Z(n2153) );
  XOR \b/SBOX[5].sbox/U117  ( .A(\b/SBOX[5].sbox/t[3] ), .B(
        \b/SBOX[5].sbox/t[8] ), .Z(n2154) );
  XOR \b/SBOX[5].sbox/U116  ( .A(n2156), .B(n2155), .Z(\b/SBOX[5].sbox/t[41] )
         );
  XOR \b/SBOX[5].sbox/U115  ( .A(n2200), .B(n2157), .Z(n2155) );
  XOR \b/SBOX[5].sbox/U114  ( .A(\b/SBOX[5].sbox/t[32] ), .B(msg[47]), .Z(
        n2156) );
  XOR \b/SBOX[5].sbox/U113  ( .A(\b/SBOX[5].sbox/t[5] ), .B(
        \b/SBOX[5].sbox/t[10] ), .Z(n2157) );
  XOR \b/SBOX[5].sbox/U112  ( .A(\b/SBOX[5].sbox/t[2] ), .B(msg[46]), .Z(n2201) );
  XOR \b/SBOX[5].sbox/U111  ( .A(n2159), .B(n2158), .Z(\b/SBOX[5].sbox/t[45] )
         );
  XOR \b/SBOX[5].sbox/U110  ( .A(n2201), .B(n2160), .Z(n2158) );
  XOR \b/SBOX[5].sbox/U109  ( .A(msg[44]), .B(n2200), .Z(n2159) );
  XOR \b/SBOX[5].sbox/U108  ( .A(\b/SBOX[5].sbox/t[7] ), .B(
        \b/SBOX[5].sbox/t[28] ), .Z(n2160) );
  XOR \b/SBOX[5].sbox/U107  ( .A(n2201), .B(n2161), .Z(n2206) );
  XOR \b/SBOX[5].sbox/U106  ( .A(\b/SBOX[5].sbox/t[5] ), .B(msg[44]), .Z(n2161) );
  XOR \b/SBOX[5].sbox/U105  ( .A(msg[47]), .B(n2162), .Z(n2202) );
  XOR \b/SBOX[5].sbox/U104  ( .A(\b/SBOX[5].sbox/t[7] ), .B(
        \b/SBOX[5].sbox/t[10] ), .Z(n2162) );
  XOR \b/SBOX[5].sbox/U103  ( .A(n2164), .B(n2163), .Z(\b/SBOX[5].sbox/t[42] )
         );
  XOR \b/SBOX[5].sbox/U102  ( .A(n2206), .B(n2202), .Z(n2163) );
  XOR \b/SBOX[5].sbox/U101  ( .A(\b/SBOX[5].sbox/t[28] ), .B(
        \b/SBOX[5].sbox/t[32] ), .Z(n2164) );
  XOR \b/SBOX[5].sbox/U100  ( .A(msg[41]), .B(n2165), .Z(n2204) );
  XOR \b/SBOX[5].sbox/U99  ( .A(msg[43]), .B(msg[42]), .Z(n2165) );
  XOR \b/SBOX[5].sbox/U98  ( .A(msg[45]), .B(n2204), .Z(\b/SBOX[5].sbox/y[16] ) );
  XOR \b/SBOX[5].sbox/U97  ( .A(\b/SBOX[5].sbox/y[16] ), .B(n2166), .Z(n2205)
         );
  XOR \b/SBOX[5].sbox/U96  ( .A(\b/SBOX[5].sbox/t[12] ), .B(
        \b/SBOX[5].sbox/t[15] ), .Z(n2166) );
  XOR \b/SBOX[5].sbox/U95  ( .A(n2205), .B(n2167), .Z(\b/SBOX[5].sbox/t[29] )
         );
  XOR \b/SBOX[5].sbox/U94  ( .A(\b/SBOX[5].sbox/t[28] ), .B(n2206), .Z(n2167)
         );
  XOR \b/SBOX[5].sbox/U93  ( .A(msg[40]), .B(n2168), .Z(\b/SBOX[5].sbox/y[1] )
         );
  XOR \b/SBOX[5].sbox/U92  ( .A(msg[46]), .B(msg[45]), .Z(n2168) );
  XOR \b/SBOX[5].sbox/U91  ( .A(msg[47]), .B(\b/SBOX[5].sbox/y[1] ), .Z(
        \b/SBOX[5].sbox/y[2] ) );
  XOR \b/SBOX[5].sbox/U90  ( .A(n2170), .B(n2169), .Z(\b/SBOX[5].sbox/t[25] )
         );
  XOR \b/SBOX[5].sbox/U89  ( .A(n2172), .B(n2171), .Z(n2169) );
  XOR \b/SBOX[5].sbox/U88  ( .A(msg[47]), .B(msg[45]), .Z(n2170) );
  XOR \b/SBOX[5].sbox/U87  ( .A(\b/SBOX[5].sbox/t[13] ), .B(
        \b/SBOX[5].sbox/t[15] ), .Z(n2171) );
  XOR \b/SBOX[5].sbox/U86  ( .A(\b/SBOX[5].sbox/t[3] ), .B(
        \b/SBOX[5].sbox/t[5] ), .Z(n2172) );
  XOR \b/SBOX[5].sbox/U85  ( .A(\b/SBOX[5].sbox/t[39] ), .B(
        \b/SBOX[5].sbox/t[25] ), .Z(\b/SBOX[5].sbox/t[40] ) );
  XOR \b/SBOX[5].sbox/U84  ( .A(msg[41]), .B(\b/SBOX[5].sbox/y[1] ), .Z(
        \b/SBOX[5].sbox/y[5] ) );
  XOR \b/SBOX[5].sbox/U83  ( .A(n2174), .B(n2173), .Z(\b/SBOX[5].sbox/y[15] )
         );
  XOR \b/SBOX[5].sbox/U82  ( .A(msg[43]), .B(msg[41]), .Z(n2173) );
  XOR \b/SBOX[5].sbox/U81  ( .A(msg[47]), .B(msg[44]), .Z(n2174) );
  XOR \b/SBOX[5].sbox/U80  ( .A(n2176), .B(n2175), .Z(\b/SBOX[5].sbox/t[21] )
         );
  XOR \b/SBOX[5].sbox/U79  ( .A(n2178), .B(n2177), .Z(n2175) );
  XOR \b/SBOX[5].sbox/U78  ( .A(\b/SBOX[5].sbox/y[15] ), .B(n2201), .Z(n2176)
         );
  XOR \b/SBOX[5].sbox/U77  ( .A(\b/SBOX[5].sbox/t[13] ), .B(msg[42]), .Z(n2177) );
  XOR \b/SBOX[5].sbox/U76  ( .A(\b/SBOX[5].sbox/t[3] ), .B(
        \b/SBOX[5].sbox/t[12] ), .Z(n2178) );
  XOR \b/SBOX[5].sbox/U75  ( .A(\b/SBOX[5].sbox/t[21] ), .B(n2179), .Z(
        \b/SBOX[5].sbox/t[43] ) );
  XOR \b/SBOX[5].sbox/U74  ( .A(\b/SBOX[5].sbox/t[28] ), .B(
        \b/SBOX[5].sbox/t[39] ), .Z(n2179) );
  XOR \b/SBOX[5].sbox/U73  ( .A(n2205), .B(n2202), .Z(\b/SBOX[5].sbox/t[24] )
         );
  XOR \b/SBOX[5].sbox/U72  ( .A(\b/SBOX[5].sbox/t[32] ), .B(
        \b/SBOX[5].sbox/t[24] ), .Z(\b/SBOX[5].sbox/t[33] ) );
  XOR \b/SBOX[5].sbox/U71  ( .A(msg[44]), .B(\b/SBOX[5].sbox/y[1] ), .Z(
        \b/SBOX[5].sbox/y[4] ) );
  XOR \b/SBOX[5].sbox/U70  ( .A(n2181), .B(n2180), .Z(\b/SBOX[5].sbox/t[30] )
         );
  XOR \b/SBOX[5].sbox/U69  ( .A(msg[41]), .B(n2182), .Z(n2180) );
  XOR \b/SBOX[5].sbox/U68  ( .A(\b/SBOX[5].sbox/t[13] ), .B(
        \b/SBOX[5].sbox/t[15] ), .Z(n2181) );
  XOR \b/SBOX[5].sbox/U67  ( .A(\b/SBOX[5].sbox/t[8] ), .B(
        \b/SBOX[5].sbox/t[10] ), .Z(n2182) );
  XOR \b/SBOX[5].sbox/U66  ( .A(\b/SBOX[5].sbox/t[30] ), .B(n2183), .Z(
        \b/SBOX[5].sbox/t[37] ) );
  XOR \b/SBOX[5].sbox/U65  ( .A(\b/SBOX[5].sbox/t[32] ), .B(
        \b/SBOX[5].sbox/t[36] ), .Z(n2183) );
  XOR \b/SBOX[5].sbox/U64  ( .A(msg[47]), .B(msg[42]), .Z(n2203) );
  XOR \b/SBOX[5].sbox/U63  ( .A(\b/SBOX[5].sbox/y[5] ), .B(n2203), .Z(
        \b/SBOX[5].sbox/y[3] ) );
  XOR \b/SBOX[5].sbox/U62  ( .A(n2185), .B(n2184), .Z(\b/SBOX[5].sbox/t[23] )
         );
  XOR \b/SBOX[5].sbox/U61  ( .A(n2187), .B(n2186), .Z(n2184) );
  XOR \b/SBOX[5].sbox/U60  ( .A(n2203), .B(n2188), .Z(n2185) );
  XOR \b/SBOX[5].sbox/U59  ( .A(msg[45]), .B(msg[43]), .Z(n2186) );
  XOR \b/SBOX[5].sbox/U58  ( .A(\b/SBOX[5].sbox/t[12] ), .B(
        \b/SBOX[5].sbox/t[13] ), .Z(n2187) );
  XOR \b/SBOX[5].sbox/U57  ( .A(\b/SBOX[5].sbox/t[7] ), .B(
        \b/SBOX[5].sbox/t[8] ), .Z(n2188) );
  XOR \b/SBOX[5].sbox/U56  ( .A(\b/SBOX[5].sbox/t[36] ), .B(
        \b/SBOX[5].sbox/t[23] ), .Z(\b/SBOX[5].sbox/t[44] ) );
  XOR \b/SBOX[5].sbox/U55  ( .A(n2203), .B(n2189), .Z(\b/SBOX[5].sbox/y[12] )
         );
  XOR \b/SBOX[5].sbox/U54  ( .A(msg[44]), .B(msg[41]), .Z(n2189) );
  XOR \b/SBOX[5].sbox/U53  ( .A(\b/SBOX[5].sbox/y[15] ), .B(n2190), .Z(
        \b/SBOX[5].sbox/y[10] ) );
  XOR \b/SBOX[5].sbox/U52  ( .A(msg[46]), .B(msg[45]), .Z(n2190) );
  XOR \b/SBOX[5].sbox/U51  ( .A(n2203), .B(n2191), .Z(\b/SBOX[5].sbox/y[17] )
         );
  XOR \b/SBOX[5].sbox/U50  ( .A(msg[45]), .B(msg[44]), .Z(n2191) );
  XOR \b/SBOX[5].sbox/U49  ( .A(msg[46]), .B(n2204), .Z(\b/SBOX[5].sbox/y[11] ) );
  XOR \b/SBOX[5].sbox/U48  ( .A(msg[40]), .B(\b/SBOX[5].sbox/y[11] ), .Z(
        \b/SBOX[5].sbox/y[7] ) );
  XOR \b/SBOX[5].sbox/U47  ( .A(msg[40]), .B(\b/SBOX[5].sbox/y[15] ), .Z(
        \b/SBOX[5].sbox/y[6] ) );
  XOR \b/SBOX[5].sbox/U46  ( .A(\b/SBOX[5].sbox/t[26] ), .B(
        \b/SBOX[5].sbox/t[24] ), .Z(\b/SBOX[5].sbox/t[27] ) );
  XOR \b/SBOX[5].sbox/U45  ( .A(\b/SBOX[5].sbox/t[36] ), .B(
        \b/SBOX[5].sbox/t[27] ), .Z(\b/SBOX[5].sbox/t[38] ) );
  XOR \b/SBOX[5].sbox/U44  ( .A(n2205), .B(n2192), .Z(\b/SBOX[5].sbox/t[31] )
         );
  XOR \b/SBOX[5].sbox/U43  ( .A(\b/SBOX[5].sbox/t[26] ), .B(n2206), .Z(n2192)
         );
  XOR \b/SBOX[4].sbox/U157  ( .A(\b/SBOX[4].sbox/z[12] ), .B(n2049), .Z(n2113)
         );
  XOR \b/SBOX[4].sbox/U156  ( .A(\b/SBOX[4].sbox/z[0] ), .B(
        \b/SBOX[4].sbox/z[2] ), .Z(n2049) );
  XOR \b/SBOX[4].sbox/U155  ( .A(n2051), .B(n2050), .Z(n2112) );
  XOR \b/SBOX[4].sbox/U154  ( .A(\b/SBOX[4].sbox/z[15] ), .B(
        \b/SBOX[4].sbox/z[16] ), .Z(n2050) );
  XOR \b/SBOX[4].sbox/U153  ( .A(\b/SBOX[4].sbox/z[5] ), .B(
        \b/SBOX[4].sbox/z[13] ), .Z(n2051) );
  XOR \b/SBOX[4].sbox/U152  ( .A(n2112), .B(n2052), .Z(n2126) );
  XOR \b/SBOX[4].sbox/U151  ( .A(\b/SBOX[4].sbox/z[3] ), .B(n2113), .Z(n2052)
         );
  XOR \b/SBOX[4].sbox/U150  ( .A(n2054), .B(n2053), .Z(n2127) );
  XOR \b/SBOX[4].sbox/U149  ( .A(n2112), .B(n2055), .Z(n2053) );
  XOR \b/SBOX[4].sbox/U148  ( .A(\b/SBOX[4].sbox/z[8] ), .B(
        \b/SBOX[4].sbox/z[12] ), .Z(n2054) );
  XOR \b/SBOX[4].sbox/U147  ( .A(\b/SBOX[4].sbox/z[4] ), .B(
        \b/SBOX[4].sbox/z[7] ), .Z(n2055) );
  XOR \b/SBOX[4].sbox/U146  ( .A(n2113), .B(n2056), .Z(n2115) );
  XOR \b/SBOX[4].sbox/U145  ( .A(\b/SBOX[4].sbox/z[8] ), .B(
        \b/SBOX[4].sbox/z[14] ), .Z(n2056) );
  XOR \b/SBOX[4].sbox/U144  ( .A(n2058), .B(n2057), .Z(n2128) );
  XOR \b/SBOX[4].sbox/U143  ( .A(\b/SBOX[4].sbox/z[17] ), .B(n2115), .Z(n2057)
         );
  XOR \b/SBOX[4].sbox/U142  ( .A(\b/SBOX[4].sbox/z[6] ), .B(
        \b/SBOX[4].sbox/z[15] ), .Z(n2058) );
  XOR \b/SBOX[4].sbox/U141  ( .A(\b/SBOX[4].sbox/z[9] ), .B(n2059), .Z(n2116)
         );
  XOR \b/SBOX[4].sbox/U140  ( .A(\b/SBOX[4].sbox/z[0] ), .B(
        \b/SBOX[4].sbox/z[1] ), .Z(n2059) );
  XOR \b/SBOX[4].sbox/U139  ( .A(\b/SBOX[4].sbox/z[16] ), .B(n2060), .Z(n2114)
         );
  XOR \b/SBOX[4].sbox/U138  ( .A(\b/SBOX[4].sbox/z[10] ), .B(
        \b/SBOX[4].sbox/z[15] ), .Z(n2060) );
  XOR \b/SBOX[4].sbox/U137  ( .A(n2062), .B(n2061), .Z(n2129) );
  XOR \b/SBOX[4].sbox/U136  ( .A(n2116), .B(n2114), .Z(n2061) );
  XOR \b/SBOX[4].sbox/U135  ( .A(\b/SBOX[4].sbox/z[6] ), .B(
        \b/SBOX[4].sbox/z[7] ), .Z(n2062) );
  XOR \b/SBOX[4].sbox/U134  ( .A(\b/SBOX[4].sbox/z[4] ), .B(n2114), .Z(n2117)
         );
  XOR \b/SBOX[4].sbox/U133  ( .A(n2117), .B(n2063), .Z(n2118) );
  XOR \b/SBOX[4].sbox/U132  ( .A(\b/SBOX[4].sbox/z[3] ), .B(
        \b/SBOX[4].sbox/z[7] ), .Z(n2063) );
  XOR \b/SBOX[4].sbox/U131  ( .A(n2115), .B(n2064), .Z(shift_row_out[34]) );
  XOR \b/SBOX[4].sbox/U130  ( .A(\b/SBOX[4].sbox/z[11] ), .B(n2118), .Z(n2064)
         );
  XOR \b/SBOX[4].sbox/U129  ( .A(n2066), .B(n2065), .Z(shift_row_out[35]) );
  XOR \b/SBOX[4].sbox/U128  ( .A(n2117), .B(n2067), .Z(n2065) );
  XOR \b/SBOX[4].sbox/U127  ( .A(\b/SBOX[4].sbox/z[5] ), .B(
        \b/SBOX[4].sbox/z[9] ), .Z(n2066) );
  XOR \b/SBOX[4].sbox/U126  ( .A(\b/SBOX[4].sbox/z[1] ), .B(
        \b/SBOX[4].sbox/z[2] ), .Z(n2067) );
  XOR \b/SBOX[4].sbox/U125  ( .A(n2116), .B(n2068), .Z(shift_row_out[36]) );
  XOR \b/SBOX[4].sbox/U124  ( .A(\b/SBOX[4].sbox/z[3] ), .B(n2117), .Z(n2068)
         );
  XOR \b/SBOX[4].sbox/U123  ( .A(n2118), .B(n2069), .Z(shift_row_out[39]) );
  XOR \b/SBOX[4].sbox/U122  ( .A(\b/SBOX[4].sbox/z[6] ), .B(
        \b/SBOX[4].sbox/z[9] ), .Z(n2069) );
  XOR \b/SBOX[4].sbox/U121  ( .A(n2071), .B(n2070), .Z(n2119) );
  XOR \b/SBOX[4].sbox/U120  ( .A(n2073), .B(n2072), .Z(n2070) );
  XOR \b/SBOX[4].sbox/U119  ( .A(msg[37]), .B(msg[33]), .Z(n2071) );
  XOR \b/SBOX[4].sbox/U118  ( .A(\b/SBOX[4].sbox/t[36] ), .B(
        \b/SBOX[4].sbox/t[39] ), .Z(n2072) );
  XOR \b/SBOX[4].sbox/U117  ( .A(\b/SBOX[4].sbox/t[3] ), .B(
        \b/SBOX[4].sbox/t[8] ), .Z(n2073) );
  XOR \b/SBOX[4].sbox/U116  ( .A(n2075), .B(n2074), .Z(\b/SBOX[4].sbox/t[41] )
         );
  XOR \b/SBOX[4].sbox/U115  ( .A(n2119), .B(n2076), .Z(n2074) );
  XOR \b/SBOX[4].sbox/U114  ( .A(\b/SBOX[4].sbox/t[32] ), .B(msg[39]), .Z(
        n2075) );
  XOR \b/SBOX[4].sbox/U113  ( .A(\b/SBOX[4].sbox/t[5] ), .B(
        \b/SBOX[4].sbox/t[10] ), .Z(n2076) );
  XOR \b/SBOX[4].sbox/U112  ( .A(\b/SBOX[4].sbox/t[2] ), .B(msg[38]), .Z(n2120) );
  XOR \b/SBOX[4].sbox/U111  ( .A(n2078), .B(n2077), .Z(\b/SBOX[4].sbox/t[45] )
         );
  XOR \b/SBOX[4].sbox/U110  ( .A(n2120), .B(n2079), .Z(n2077) );
  XOR \b/SBOX[4].sbox/U109  ( .A(msg[36]), .B(n2119), .Z(n2078) );
  XOR \b/SBOX[4].sbox/U108  ( .A(\b/SBOX[4].sbox/t[7] ), .B(
        \b/SBOX[4].sbox/t[28] ), .Z(n2079) );
  XOR \b/SBOX[4].sbox/U107  ( .A(n2120), .B(n2080), .Z(n2125) );
  XOR \b/SBOX[4].sbox/U106  ( .A(\b/SBOX[4].sbox/t[5] ), .B(msg[36]), .Z(n2080) );
  XOR \b/SBOX[4].sbox/U105  ( .A(msg[39]), .B(n2081), .Z(n2121) );
  XOR \b/SBOX[4].sbox/U104  ( .A(\b/SBOX[4].sbox/t[7] ), .B(
        \b/SBOX[4].sbox/t[10] ), .Z(n2081) );
  XOR \b/SBOX[4].sbox/U103  ( .A(n2083), .B(n2082), .Z(\b/SBOX[4].sbox/t[42] )
         );
  XOR \b/SBOX[4].sbox/U102  ( .A(n2125), .B(n2121), .Z(n2082) );
  XOR \b/SBOX[4].sbox/U101  ( .A(\b/SBOX[4].sbox/t[28] ), .B(
        \b/SBOX[4].sbox/t[32] ), .Z(n2083) );
  XOR \b/SBOX[4].sbox/U100  ( .A(msg[33]), .B(n2084), .Z(n2123) );
  XOR \b/SBOX[4].sbox/U99  ( .A(msg[35]), .B(msg[34]), .Z(n2084) );
  XOR \b/SBOX[4].sbox/U98  ( .A(msg[37]), .B(n2123), .Z(\b/SBOX[4].sbox/y[16] ) );
  XOR \b/SBOX[4].sbox/U97  ( .A(\b/SBOX[4].sbox/y[16] ), .B(n2085), .Z(n2124)
         );
  XOR \b/SBOX[4].sbox/U96  ( .A(\b/SBOX[4].sbox/t[12] ), .B(
        \b/SBOX[4].sbox/t[15] ), .Z(n2085) );
  XOR \b/SBOX[4].sbox/U95  ( .A(n2124), .B(n2086), .Z(\b/SBOX[4].sbox/t[29] )
         );
  XOR \b/SBOX[4].sbox/U94  ( .A(\b/SBOX[4].sbox/t[28] ), .B(n2125), .Z(n2086)
         );
  XOR \b/SBOX[4].sbox/U93  ( .A(msg[32]), .B(n2087), .Z(\b/SBOX[4].sbox/y[1] )
         );
  XOR \b/SBOX[4].sbox/U92  ( .A(msg[38]), .B(msg[37]), .Z(n2087) );
  XOR \b/SBOX[4].sbox/U91  ( .A(msg[39]), .B(\b/SBOX[4].sbox/y[1] ), .Z(
        \b/SBOX[4].sbox/y[2] ) );
  XOR \b/SBOX[4].sbox/U90  ( .A(n2089), .B(n2088), .Z(\b/SBOX[4].sbox/t[25] )
         );
  XOR \b/SBOX[4].sbox/U89  ( .A(n2091), .B(n2090), .Z(n2088) );
  XOR \b/SBOX[4].sbox/U88  ( .A(msg[39]), .B(msg[37]), .Z(n2089) );
  XOR \b/SBOX[4].sbox/U87  ( .A(\b/SBOX[4].sbox/t[13] ), .B(
        \b/SBOX[4].sbox/t[15] ), .Z(n2090) );
  XOR \b/SBOX[4].sbox/U86  ( .A(\b/SBOX[4].sbox/t[3] ), .B(
        \b/SBOX[4].sbox/t[5] ), .Z(n2091) );
  XOR \b/SBOX[4].sbox/U85  ( .A(\b/SBOX[4].sbox/t[39] ), .B(
        \b/SBOX[4].sbox/t[25] ), .Z(\b/SBOX[4].sbox/t[40] ) );
  XOR \b/SBOX[4].sbox/U84  ( .A(msg[33]), .B(\b/SBOX[4].sbox/y[1] ), .Z(
        \b/SBOX[4].sbox/y[5] ) );
  XOR \b/SBOX[4].sbox/U83  ( .A(n2093), .B(n2092), .Z(\b/SBOX[4].sbox/y[15] )
         );
  XOR \b/SBOX[4].sbox/U82  ( .A(msg[35]), .B(msg[33]), .Z(n2092) );
  XOR \b/SBOX[4].sbox/U81  ( .A(msg[39]), .B(msg[36]), .Z(n2093) );
  XOR \b/SBOX[4].sbox/U80  ( .A(n2095), .B(n2094), .Z(\b/SBOX[4].sbox/t[21] )
         );
  XOR \b/SBOX[4].sbox/U79  ( .A(n2097), .B(n2096), .Z(n2094) );
  XOR \b/SBOX[4].sbox/U78  ( .A(\b/SBOX[4].sbox/y[15] ), .B(n2120), .Z(n2095)
         );
  XOR \b/SBOX[4].sbox/U77  ( .A(\b/SBOX[4].sbox/t[13] ), .B(msg[34]), .Z(n2096) );
  XOR \b/SBOX[4].sbox/U76  ( .A(\b/SBOX[4].sbox/t[3] ), .B(
        \b/SBOX[4].sbox/t[12] ), .Z(n2097) );
  XOR \b/SBOX[4].sbox/U75  ( .A(\b/SBOX[4].sbox/t[21] ), .B(n2098), .Z(
        \b/SBOX[4].sbox/t[43] ) );
  XOR \b/SBOX[4].sbox/U74  ( .A(\b/SBOX[4].sbox/t[28] ), .B(
        \b/SBOX[4].sbox/t[39] ), .Z(n2098) );
  XOR \b/SBOX[4].sbox/U73  ( .A(n2124), .B(n2121), .Z(\b/SBOX[4].sbox/t[24] )
         );
  XOR \b/SBOX[4].sbox/U72  ( .A(\b/SBOX[4].sbox/t[32] ), .B(
        \b/SBOX[4].sbox/t[24] ), .Z(\b/SBOX[4].sbox/t[33] ) );
  XOR \b/SBOX[4].sbox/U71  ( .A(msg[36]), .B(\b/SBOX[4].sbox/y[1] ), .Z(
        \b/SBOX[4].sbox/y[4] ) );
  XOR \b/SBOX[4].sbox/U70  ( .A(n2100), .B(n2099), .Z(\b/SBOX[4].sbox/t[30] )
         );
  XOR \b/SBOX[4].sbox/U69  ( .A(msg[33]), .B(n2101), .Z(n2099) );
  XOR \b/SBOX[4].sbox/U68  ( .A(\b/SBOX[4].sbox/t[13] ), .B(
        \b/SBOX[4].sbox/t[15] ), .Z(n2100) );
  XOR \b/SBOX[4].sbox/U67  ( .A(\b/SBOX[4].sbox/t[8] ), .B(
        \b/SBOX[4].sbox/t[10] ), .Z(n2101) );
  XOR \b/SBOX[4].sbox/U66  ( .A(\b/SBOX[4].sbox/t[30] ), .B(n2102), .Z(
        \b/SBOX[4].sbox/t[37] ) );
  XOR \b/SBOX[4].sbox/U65  ( .A(\b/SBOX[4].sbox/t[32] ), .B(
        \b/SBOX[4].sbox/t[36] ), .Z(n2102) );
  XOR \b/SBOX[4].sbox/U64  ( .A(msg[39]), .B(msg[34]), .Z(n2122) );
  XOR \b/SBOX[4].sbox/U63  ( .A(\b/SBOX[4].sbox/y[5] ), .B(n2122), .Z(
        \b/SBOX[4].sbox/y[3] ) );
  XOR \b/SBOX[4].sbox/U62  ( .A(n2104), .B(n2103), .Z(\b/SBOX[4].sbox/t[23] )
         );
  XOR \b/SBOX[4].sbox/U61  ( .A(n2106), .B(n2105), .Z(n2103) );
  XOR \b/SBOX[4].sbox/U60  ( .A(n2122), .B(n2107), .Z(n2104) );
  XOR \b/SBOX[4].sbox/U59  ( .A(msg[37]), .B(msg[35]), .Z(n2105) );
  XOR \b/SBOX[4].sbox/U58  ( .A(\b/SBOX[4].sbox/t[12] ), .B(
        \b/SBOX[4].sbox/t[13] ), .Z(n2106) );
  XOR \b/SBOX[4].sbox/U57  ( .A(\b/SBOX[4].sbox/t[7] ), .B(
        \b/SBOX[4].sbox/t[8] ), .Z(n2107) );
  XOR \b/SBOX[4].sbox/U56  ( .A(\b/SBOX[4].sbox/t[36] ), .B(
        \b/SBOX[4].sbox/t[23] ), .Z(\b/SBOX[4].sbox/t[44] ) );
  XOR \b/SBOX[4].sbox/U55  ( .A(n2122), .B(n2108), .Z(\b/SBOX[4].sbox/y[12] )
         );
  XOR \b/SBOX[4].sbox/U54  ( .A(msg[36]), .B(msg[33]), .Z(n2108) );
  XOR \b/SBOX[4].sbox/U53  ( .A(\b/SBOX[4].sbox/y[15] ), .B(n2109), .Z(
        \b/SBOX[4].sbox/y[10] ) );
  XOR \b/SBOX[4].sbox/U52  ( .A(msg[38]), .B(msg[37]), .Z(n2109) );
  XOR \b/SBOX[4].sbox/U51  ( .A(n2122), .B(n2110), .Z(\b/SBOX[4].sbox/y[17] )
         );
  XOR \b/SBOX[4].sbox/U50  ( .A(msg[37]), .B(msg[36]), .Z(n2110) );
  XOR \b/SBOX[4].sbox/U49  ( .A(msg[38]), .B(n2123), .Z(\b/SBOX[4].sbox/y[11] ) );
  XOR \b/SBOX[4].sbox/U48  ( .A(msg[32]), .B(\b/SBOX[4].sbox/y[11] ), .Z(
        \b/SBOX[4].sbox/y[7] ) );
  XOR \b/SBOX[4].sbox/U47  ( .A(msg[32]), .B(\b/SBOX[4].sbox/y[15] ), .Z(
        \b/SBOX[4].sbox/y[6] ) );
  XOR \b/SBOX[4].sbox/U46  ( .A(\b/SBOX[4].sbox/t[26] ), .B(
        \b/SBOX[4].sbox/t[24] ), .Z(\b/SBOX[4].sbox/t[27] ) );
  XOR \b/SBOX[4].sbox/U45  ( .A(\b/SBOX[4].sbox/t[36] ), .B(
        \b/SBOX[4].sbox/t[27] ), .Z(\b/SBOX[4].sbox/t[38] ) );
  XOR \b/SBOX[4].sbox/U44  ( .A(n2124), .B(n2111), .Z(\b/SBOX[4].sbox/t[31] )
         );
  XOR \b/SBOX[4].sbox/U43  ( .A(\b/SBOX[4].sbox/t[26] ), .B(n2125), .Z(n2111)
         );
  XOR \b/SBOX[3].sbox/U157  ( .A(\b/SBOX[3].sbox/z[12] ), .B(n1968), .Z(n2032)
         );
  XOR \b/SBOX[3].sbox/U156  ( .A(\b/SBOX[3].sbox/z[0] ), .B(
        \b/SBOX[3].sbox/z[2] ), .Z(n1968) );
  XOR \b/SBOX[3].sbox/U155  ( .A(n1970), .B(n1969), .Z(n2031) );
  XOR \b/SBOX[3].sbox/U154  ( .A(\b/SBOX[3].sbox/z[15] ), .B(
        \b/SBOX[3].sbox/z[16] ), .Z(n1969) );
  XOR \b/SBOX[3].sbox/U153  ( .A(\b/SBOX[3].sbox/z[5] ), .B(
        \b/SBOX[3].sbox/z[13] ), .Z(n1970) );
  XOR \b/SBOX[3].sbox/U152  ( .A(n2031), .B(n1971), .Z(n2045) );
  XOR \b/SBOX[3].sbox/U151  ( .A(\b/SBOX[3].sbox/z[3] ), .B(n2032), .Z(n1971)
         );
  XOR \b/SBOX[3].sbox/U150  ( .A(n1973), .B(n1972), .Z(n2046) );
  XOR \b/SBOX[3].sbox/U149  ( .A(n2031), .B(n1974), .Z(n1972) );
  XOR \b/SBOX[3].sbox/U148  ( .A(\b/SBOX[3].sbox/z[8] ), .B(
        \b/SBOX[3].sbox/z[12] ), .Z(n1973) );
  XOR \b/SBOX[3].sbox/U147  ( .A(\b/SBOX[3].sbox/z[4] ), .B(
        \b/SBOX[3].sbox/z[7] ), .Z(n1974) );
  XOR \b/SBOX[3].sbox/U146  ( .A(n2032), .B(n1975), .Z(n2034) );
  XOR \b/SBOX[3].sbox/U145  ( .A(\b/SBOX[3].sbox/z[8] ), .B(
        \b/SBOX[3].sbox/z[14] ), .Z(n1975) );
  XOR \b/SBOX[3].sbox/U144  ( .A(n1977), .B(n1976), .Z(n2047) );
  XOR \b/SBOX[3].sbox/U143  ( .A(\b/SBOX[3].sbox/z[17] ), .B(n2034), .Z(n1976)
         );
  XOR \b/SBOX[3].sbox/U142  ( .A(\b/SBOX[3].sbox/z[6] ), .B(
        \b/SBOX[3].sbox/z[15] ), .Z(n1977) );
  XOR \b/SBOX[3].sbox/U141  ( .A(\b/SBOX[3].sbox/z[9] ), .B(n1978), .Z(n2035)
         );
  XOR \b/SBOX[3].sbox/U140  ( .A(\b/SBOX[3].sbox/z[0] ), .B(
        \b/SBOX[3].sbox/z[1] ), .Z(n1978) );
  XOR \b/SBOX[3].sbox/U139  ( .A(\b/SBOX[3].sbox/z[16] ), .B(n1979), .Z(n2033)
         );
  XOR \b/SBOX[3].sbox/U138  ( .A(\b/SBOX[3].sbox/z[10] ), .B(
        \b/SBOX[3].sbox/z[15] ), .Z(n1979) );
  XOR \b/SBOX[3].sbox/U137  ( .A(n1981), .B(n1980), .Z(n2048) );
  XOR \b/SBOX[3].sbox/U136  ( .A(n2035), .B(n2033), .Z(n1980) );
  XOR \b/SBOX[3].sbox/U135  ( .A(\b/SBOX[3].sbox/z[6] ), .B(
        \b/SBOX[3].sbox/z[7] ), .Z(n1981) );
  XOR \b/SBOX[3].sbox/U134  ( .A(\b/SBOX[3].sbox/z[4] ), .B(n2033), .Z(n2036)
         );
  XOR \b/SBOX[3].sbox/U133  ( .A(n2036), .B(n1982), .Z(n2037) );
  XOR \b/SBOX[3].sbox/U132  ( .A(\b/SBOX[3].sbox/z[3] ), .B(
        \b/SBOX[3].sbox/z[7] ), .Z(n1982) );
  XOR \b/SBOX[3].sbox/U131  ( .A(n2034), .B(n1983), .Z(shift_row_out[58]) );
  XOR \b/SBOX[3].sbox/U130  ( .A(\b/SBOX[3].sbox/z[11] ), .B(n2037), .Z(n1983)
         );
  XOR \b/SBOX[3].sbox/U129  ( .A(n1985), .B(n1984), .Z(shift_row_out[59]) );
  XOR \b/SBOX[3].sbox/U128  ( .A(n2036), .B(n1986), .Z(n1984) );
  XOR \b/SBOX[3].sbox/U127  ( .A(\b/SBOX[3].sbox/z[5] ), .B(
        \b/SBOX[3].sbox/z[9] ), .Z(n1985) );
  XOR \b/SBOX[3].sbox/U126  ( .A(\b/SBOX[3].sbox/z[1] ), .B(
        \b/SBOX[3].sbox/z[2] ), .Z(n1986) );
  XOR \b/SBOX[3].sbox/U125  ( .A(n2035), .B(n1987), .Z(shift_row_out[60]) );
  XOR \b/SBOX[3].sbox/U124  ( .A(\b/SBOX[3].sbox/z[3] ), .B(n2036), .Z(n1987)
         );
  XOR \b/SBOX[3].sbox/U123  ( .A(n2037), .B(n1988), .Z(shift_row_out[63]) );
  XOR \b/SBOX[3].sbox/U122  ( .A(\b/SBOX[3].sbox/z[6] ), .B(
        \b/SBOX[3].sbox/z[9] ), .Z(n1988) );
  XOR \b/SBOX[3].sbox/U121  ( .A(n1990), .B(n1989), .Z(n2038) );
  XOR \b/SBOX[3].sbox/U120  ( .A(n1992), .B(n1991), .Z(n1989) );
  XOR \b/SBOX[3].sbox/U119  ( .A(msg[29]), .B(msg[25]), .Z(n1990) );
  XOR \b/SBOX[3].sbox/U118  ( .A(\b/SBOX[3].sbox/t[36] ), .B(
        \b/SBOX[3].sbox/t[39] ), .Z(n1991) );
  XOR \b/SBOX[3].sbox/U117  ( .A(\b/SBOX[3].sbox/t[3] ), .B(
        \b/SBOX[3].sbox/t[8] ), .Z(n1992) );
  XOR \b/SBOX[3].sbox/U116  ( .A(n1994), .B(n1993), .Z(\b/SBOX[3].sbox/t[41] )
         );
  XOR \b/SBOX[3].sbox/U115  ( .A(n2038), .B(n1995), .Z(n1993) );
  XOR \b/SBOX[3].sbox/U114  ( .A(\b/SBOX[3].sbox/t[32] ), .B(msg[31]), .Z(
        n1994) );
  XOR \b/SBOX[3].sbox/U113  ( .A(\b/SBOX[3].sbox/t[5] ), .B(
        \b/SBOX[3].sbox/t[10] ), .Z(n1995) );
  XOR \b/SBOX[3].sbox/U112  ( .A(\b/SBOX[3].sbox/t[2] ), .B(msg[30]), .Z(n2039) );
  XOR \b/SBOX[3].sbox/U111  ( .A(n1997), .B(n1996), .Z(\b/SBOX[3].sbox/t[45] )
         );
  XOR \b/SBOX[3].sbox/U110  ( .A(n2039), .B(n1998), .Z(n1996) );
  XOR \b/SBOX[3].sbox/U109  ( .A(msg[28]), .B(n2038), .Z(n1997) );
  XOR \b/SBOX[3].sbox/U108  ( .A(\b/SBOX[3].sbox/t[7] ), .B(
        \b/SBOX[3].sbox/t[28] ), .Z(n1998) );
  XOR \b/SBOX[3].sbox/U107  ( .A(n2039), .B(n1999), .Z(n2044) );
  XOR \b/SBOX[3].sbox/U106  ( .A(\b/SBOX[3].sbox/t[5] ), .B(msg[28]), .Z(n1999) );
  XOR \b/SBOX[3].sbox/U105  ( .A(msg[31]), .B(n2000), .Z(n2040) );
  XOR \b/SBOX[3].sbox/U104  ( .A(\b/SBOX[3].sbox/t[7] ), .B(
        \b/SBOX[3].sbox/t[10] ), .Z(n2000) );
  XOR \b/SBOX[3].sbox/U103  ( .A(n2002), .B(n2001), .Z(\b/SBOX[3].sbox/t[42] )
         );
  XOR \b/SBOX[3].sbox/U102  ( .A(n2044), .B(n2040), .Z(n2001) );
  XOR \b/SBOX[3].sbox/U101  ( .A(\b/SBOX[3].sbox/t[28] ), .B(
        \b/SBOX[3].sbox/t[32] ), .Z(n2002) );
  XOR \b/SBOX[3].sbox/U100  ( .A(msg[25]), .B(n2003), .Z(n2042) );
  XOR \b/SBOX[3].sbox/U99  ( .A(msg[27]), .B(msg[26]), .Z(n2003) );
  XOR \b/SBOX[3].sbox/U98  ( .A(msg[29]), .B(n2042), .Z(\b/SBOX[3].sbox/y[16] ) );
  XOR \b/SBOX[3].sbox/U97  ( .A(\b/SBOX[3].sbox/y[16] ), .B(n2004), .Z(n2043)
         );
  XOR \b/SBOX[3].sbox/U96  ( .A(\b/SBOX[3].sbox/t[12] ), .B(
        \b/SBOX[3].sbox/t[15] ), .Z(n2004) );
  XOR \b/SBOX[3].sbox/U95  ( .A(n2043), .B(n2005), .Z(\b/SBOX[3].sbox/t[29] )
         );
  XOR \b/SBOX[3].sbox/U94  ( .A(\b/SBOX[3].sbox/t[28] ), .B(n2044), .Z(n2005)
         );
  XOR \b/SBOX[3].sbox/U93  ( .A(msg[24]), .B(n2006), .Z(\b/SBOX[3].sbox/y[1] )
         );
  XOR \b/SBOX[3].sbox/U92  ( .A(msg[30]), .B(msg[29]), .Z(n2006) );
  XOR \b/SBOX[3].sbox/U91  ( .A(msg[31]), .B(\b/SBOX[3].sbox/y[1] ), .Z(
        \b/SBOX[3].sbox/y[2] ) );
  XOR \b/SBOX[3].sbox/U90  ( .A(n2008), .B(n2007), .Z(\b/SBOX[3].sbox/t[25] )
         );
  XOR \b/SBOX[3].sbox/U89  ( .A(n2010), .B(n2009), .Z(n2007) );
  XOR \b/SBOX[3].sbox/U88  ( .A(msg[31]), .B(msg[29]), .Z(n2008) );
  XOR \b/SBOX[3].sbox/U87  ( .A(\b/SBOX[3].sbox/t[13] ), .B(
        \b/SBOX[3].sbox/t[15] ), .Z(n2009) );
  XOR \b/SBOX[3].sbox/U86  ( .A(\b/SBOX[3].sbox/t[3] ), .B(
        \b/SBOX[3].sbox/t[5] ), .Z(n2010) );
  XOR \b/SBOX[3].sbox/U85  ( .A(\b/SBOX[3].sbox/t[39] ), .B(
        \b/SBOX[3].sbox/t[25] ), .Z(\b/SBOX[3].sbox/t[40] ) );
  XOR \b/SBOX[3].sbox/U84  ( .A(msg[25]), .B(\b/SBOX[3].sbox/y[1] ), .Z(
        \b/SBOX[3].sbox/y[5] ) );
  XOR \b/SBOX[3].sbox/U83  ( .A(n2012), .B(n2011), .Z(\b/SBOX[3].sbox/y[15] )
         );
  XOR \b/SBOX[3].sbox/U82  ( .A(msg[27]), .B(msg[25]), .Z(n2011) );
  XOR \b/SBOX[3].sbox/U81  ( .A(msg[31]), .B(msg[28]), .Z(n2012) );
  XOR \b/SBOX[3].sbox/U80  ( .A(n2014), .B(n2013), .Z(\b/SBOX[3].sbox/t[21] )
         );
  XOR \b/SBOX[3].sbox/U79  ( .A(n2016), .B(n2015), .Z(n2013) );
  XOR \b/SBOX[3].sbox/U78  ( .A(\b/SBOX[3].sbox/y[15] ), .B(n2039), .Z(n2014)
         );
  XOR \b/SBOX[3].sbox/U77  ( .A(\b/SBOX[3].sbox/t[13] ), .B(msg[26]), .Z(n2015) );
  XOR \b/SBOX[3].sbox/U76  ( .A(\b/SBOX[3].sbox/t[3] ), .B(
        \b/SBOX[3].sbox/t[12] ), .Z(n2016) );
  XOR \b/SBOX[3].sbox/U75  ( .A(\b/SBOX[3].sbox/t[21] ), .B(n2017), .Z(
        \b/SBOX[3].sbox/t[43] ) );
  XOR \b/SBOX[3].sbox/U74  ( .A(\b/SBOX[3].sbox/t[28] ), .B(
        \b/SBOX[3].sbox/t[39] ), .Z(n2017) );
  XOR \b/SBOX[3].sbox/U73  ( .A(n2043), .B(n2040), .Z(\b/SBOX[3].sbox/t[24] )
         );
  XOR \b/SBOX[3].sbox/U72  ( .A(\b/SBOX[3].sbox/t[32] ), .B(
        \b/SBOX[3].sbox/t[24] ), .Z(\b/SBOX[3].sbox/t[33] ) );
  XOR \b/SBOX[3].sbox/U71  ( .A(msg[28]), .B(\b/SBOX[3].sbox/y[1] ), .Z(
        \b/SBOX[3].sbox/y[4] ) );
  XOR \b/SBOX[3].sbox/U70  ( .A(n2019), .B(n2018), .Z(\b/SBOX[3].sbox/t[30] )
         );
  XOR \b/SBOX[3].sbox/U69  ( .A(msg[25]), .B(n2020), .Z(n2018) );
  XOR \b/SBOX[3].sbox/U68  ( .A(\b/SBOX[3].sbox/t[13] ), .B(
        \b/SBOX[3].sbox/t[15] ), .Z(n2019) );
  XOR \b/SBOX[3].sbox/U67  ( .A(\b/SBOX[3].sbox/t[8] ), .B(
        \b/SBOX[3].sbox/t[10] ), .Z(n2020) );
  XOR \b/SBOX[3].sbox/U66  ( .A(\b/SBOX[3].sbox/t[30] ), .B(n2021), .Z(
        \b/SBOX[3].sbox/t[37] ) );
  XOR \b/SBOX[3].sbox/U65  ( .A(\b/SBOX[3].sbox/t[32] ), .B(
        \b/SBOX[3].sbox/t[36] ), .Z(n2021) );
  XOR \b/SBOX[3].sbox/U64  ( .A(msg[31]), .B(msg[26]), .Z(n2041) );
  XOR \b/SBOX[3].sbox/U63  ( .A(\b/SBOX[3].sbox/y[5] ), .B(n2041), .Z(
        \b/SBOX[3].sbox/y[3] ) );
  XOR \b/SBOX[3].sbox/U62  ( .A(n2023), .B(n2022), .Z(\b/SBOX[3].sbox/t[23] )
         );
  XOR \b/SBOX[3].sbox/U61  ( .A(n2025), .B(n2024), .Z(n2022) );
  XOR \b/SBOX[3].sbox/U60  ( .A(n2041), .B(n2026), .Z(n2023) );
  XOR \b/SBOX[3].sbox/U59  ( .A(msg[29]), .B(msg[27]), .Z(n2024) );
  XOR \b/SBOX[3].sbox/U58  ( .A(\b/SBOX[3].sbox/t[12] ), .B(
        \b/SBOX[3].sbox/t[13] ), .Z(n2025) );
  XOR \b/SBOX[3].sbox/U57  ( .A(\b/SBOX[3].sbox/t[7] ), .B(
        \b/SBOX[3].sbox/t[8] ), .Z(n2026) );
  XOR \b/SBOX[3].sbox/U56  ( .A(\b/SBOX[3].sbox/t[36] ), .B(
        \b/SBOX[3].sbox/t[23] ), .Z(\b/SBOX[3].sbox/t[44] ) );
  XOR \b/SBOX[3].sbox/U55  ( .A(n2041), .B(n2027), .Z(\b/SBOX[3].sbox/y[12] )
         );
  XOR \b/SBOX[3].sbox/U54  ( .A(msg[28]), .B(msg[25]), .Z(n2027) );
  XOR \b/SBOX[3].sbox/U53  ( .A(\b/SBOX[3].sbox/y[15] ), .B(n2028), .Z(
        \b/SBOX[3].sbox/y[10] ) );
  XOR \b/SBOX[3].sbox/U52  ( .A(msg[30]), .B(msg[29]), .Z(n2028) );
  XOR \b/SBOX[3].sbox/U51  ( .A(n2041), .B(n2029), .Z(\b/SBOX[3].sbox/y[17] )
         );
  XOR \b/SBOX[3].sbox/U50  ( .A(msg[29]), .B(msg[28]), .Z(n2029) );
  XOR \b/SBOX[3].sbox/U49  ( .A(msg[30]), .B(n2042), .Z(\b/SBOX[3].sbox/y[11] ) );
  XOR \b/SBOX[3].sbox/U48  ( .A(msg[24]), .B(\b/SBOX[3].sbox/y[11] ), .Z(
        \b/SBOX[3].sbox/y[7] ) );
  XOR \b/SBOX[3].sbox/U47  ( .A(msg[24]), .B(\b/SBOX[3].sbox/y[15] ), .Z(
        \b/SBOX[3].sbox/y[6] ) );
  XOR \b/SBOX[3].sbox/U46  ( .A(\b/SBOX[3].sbox/t[26] ), .B(
        \b/SBOX[3].sbox/t[24] ), .Z(\b/SBOX[3].sbox/t[27] ) );
  XOR \b/SBOX[3].sbox/U45  ( .A(\b/SBOX[3].sbox/t[36] ), .B(
        \b/SBOX[3].sbox/t[27] ), .Z(\b/SBOX[3].sbox/t[38] ) );
  XOR \b/SBOX[3].sbox/U44  ( .A(n2043), .B(n2030), .Z(\b/SBOX[3].sbox/t[31] )
         );
  XOR \b/SBOX[3].sbox/U43  ( .A(\b/SBOX[3].sbox/t[26] ), .B(n2044), .Z(n2030)
         );
  XOR \b/SBOX[2].sbox/U157  ( .A(\b/SBOX[2].sbox/z[12] ), .B(n1887), .Z(n1951)
         );
  XOR \b/SBOX[2].sbox/U156  ( .A(\b/SBOX[2].sbox/z[0] ), .B(
        \b/SBOX[2].sbox/z[2] ), .Z(n1887) );
  XOR \b/SBOX[2].sbox/U155  ( .A(n1889), .B(n1888), .Z(n1950) );
  XOR \b/SBOX[2].sbox/U154  ( .A(\b/SBOX[2].sbox/z[15] ), .B(
        \b/SBOX[2].sbox/z[16] ), .Z(n1888) );
  XOR \b/SBOX[2].sbox/U153  ( .A(\b/SBOX[2].sbox/z[5] ), .B(
        \b/SBOX[2].sbox/z[13] ), .Z(n1889) );
  XOR \b/SBOX[2].sbox/U152  ( .A(n1950), .B(n1890), .Z(n1964) );
  XOR \b/SBOX[2].sbox/U151  ( .A(\b/SBOX[2].sbox/z[3] ), .B(n1951), .Z(n1890)
         );
  XOR \b/SBOX[2].sbox/U150  ( .A(n1892), .B(n1891), .Z(n1965) );
  XOR \b/SBOX[2].sbox/U149  ( .A(n1950), .B(n1893), .Z(n1891) );
  XOR \b/SBOX[2].sbox/U148  ( .A(\b/SBOX[2].sbox/z[8] ), .B(
        \b/SBOX[2].sbox/z[12] ), .Z(n1892) );
  XOR \b/SBOX[2].sbox/U147  ( .A(\b/SBOX[2].sbox/z[4] ), .B(
        \b/SBOX[2].sbox/z[7] ), .Z(n1893) );
  XOR \b/SBOX[2].sbox/U146  ( .A(n1951), .B(n1894), .Z(n1953) );
  XOR \b/SBOX[2].sbox/U145  ( .A(\b/SBOX[2].sbox/z[8] ), .B(
        \b/SBOX[2].sbox/z[14] ), .Z(n1894) );
  XOR \b/SBOX[2].sbox/U144  ( .A(n1896), .B(n1895), .Z(n1966) );
  XOR \b/SBOX[2].sbox/U143  ( .A(\b/SBOX[2].sbox/z[17] ), .B(n1953), .Z(n1895)
         );
  XOR \b/SBOX[2].sbox/U142  ( .A(\b/SBOX[2].sbox/z[6] ), .B(
        \b/SBOX[2].sbox/z[15] ), .Z(n1896) );
  XOR \b/SBOX[2].sbox/U141  ( .A(\b/SBOX[2].sbox/z[9] ), .B(n1897), .Z(n1954)
         );
  XOR \b/SBOX[2].sbox/U140  ( .A(\b/SBOX[2].sbox/z[0] ), .B(
        \b/SBOX[2].sbox/z[1] ), .Z(n1897) );
  XOR \b/SBOX[2].sbox/U139  ( .A(\b/SBOX[2].sbox/z[16] ), .B(n1898), .Z(n1952)
         );
  XOR \b/SBOX[2].sbox/U138  ( .A(\b/SBOX[2].sbox/z[10] ), .B(
        \b/SBOX[2].sbox/z[15] ), .Z(n1898) );
  XOR \b/SBOX[2].sbox/U137  ( .A(n1900), .B(n1899), .Z(n1967) );
  XOR \b/SBOX[2].sbox/U136  ( .A(n1954), .B(n1952), .Z(n1899) );
  XOR \b/SBOX[2].sbox/U135  ( .A(\b/SBOX[2].sbox/z[6] ), .B(
        \b/SBOX[2].sbox/z[7] ), .Z(n1900) );
  XOR \b/SBOX[2].sbox/U134  ( .A(\b/SBOX[2].sbox/z[4] ), .B(n1952), .Z(n1955)
         );
  XOR \b/SBOX[2].sbox/U133  ( .A(n1955), .B(n1901), .Z(n1956) );
  XOR \b/SBOX[2].sbox/U132  ( .A(\b/SBOX[2].sbox/z[3] ), .B(
        \b/SBOX[2].sbox/z[7] ), .Z(n1901) );
  XOR \b/SBOX[2].sbox/U131  ( .A(n1953), .B(n1902), .Z(shift_row_out[82]) );
  XOR \b/SBOX[2].sbox/U130  ( .A(\b/SBOX[2].sbox/z[11] ), .B(n1956), .Z(n1902)
         );
  XOR \b/SBOX[2].sbox/U129  ( .A(n1904), .B(n1903), .Z(shift_row_out[83]) );
  XOR \b/SBOX[2].sbox/U128  ( .A(n1955), .B(n1905), .Z(n1903) );
  XOR \b/SBOX[2].sbox/U127  ( .A(\b/SBOX[2].sbox/z[5] ), .B(
        \b/SBOX[2].sbox/z[9] ), .Z(n1904) );
  XOR \b/SBOX[2].sbox/U126  ( .A(\b/SBOX[2].sbox/z[1] ), .B(
        \b/SBOX[2].sbox/z[2] ), .Z(n1905) );
  XOR \b/SBOX[2].sbox/U125  ( .A(n1954), .B(n1906), .Z(shift_row_out[84]) );
  XOR \b/SBOX[2].sbox/U124  ( .A(\b/SBOX[2].sbox/z[3] ), .B(n1955), .Z(n1906)
         );
  XOR \b/SBOX[2].sbox/U123  ( .A(n1956), .B(n1907), .Z(shift_row_out[87]) );
  XOR \b/SBOX[2].sbox/U122  ( .A(\b/SBOX[2].sbox/z[6] ), .B(
        \b/SBOX[2].sbox/z[9] ), .Z(n1907) );
  XOR \b/SBOX[2].sbox/U121  ( .A(n1909), .B(n1908), .Z(n1957) );
  XOR \b/SBOX[2].sbox/U120  ( .A(n1911), .B(n1910), .Z(n1908) );
  XOR \b/SBOX[2].sbox/U119  ( .A(msg[21]), .B(msg[17]), .Z(n1909) );
  XOR \b/SBOX[2].sbox/U118  ( .A(\b/SBOX[2].sbox/t[36] ), .B(
        \b/SBOX[2].sbox/t[39] ), .Z(n1910) );
  XOR \b/SBOX[2].sbox/U117  ( .A(\b/SBOX[2].sbox/t[3] ), .B(
        \b/SBOX[2].sbox/t[8] ), .Z(n1911) );
  XOR \b/SBOX[2].sbox/U116  ( .A(n1913), .B(n1912), .Z(\b/SBOX[2].sbox/t[41] )
         );
  XOR \b/SBOX[2].sbox/U115  ( .A(n1957), .B(n1914), .Z(n1912) );
  XOR \b/SBOX[2].sbox/U114  ( .A(\b/SBOX[2].sbox/t[32] ), .B(msg[23]), .Z(
        n1913) );
  XOR \b/SBOX[2].sbox/U113  ( .A(\b/SBOX[2].sbox/t[5] ), .B(
        \b/SBOX[2].sbox/t[10] ), .Z(n1914) );
  XOR \b/SBOX[2].sbox/U112  ( .A(\b/SBOX[2].sbox/t[2] ), .B(msg[22]), .Z(n1958) );
  XOR \b/SBOX[2].sbox/U111  ( .A(n1916), .B(n1915), .Z(\b/SBOX[2].sbox/t[45] )
         );
  XOR \b/SBOX[2].sbox/U110  ( .A(n1958), .B(n1917), .Z(n1915) );
  XOR \b/SBOX[2].sbox/U109  ( .A(msg[20]), .B(n1957), .Z(n1916) );
  XOR \b/SBOX[2].sbox/U108  ( .A(\b/SBOX[2].sbox/t[7] ), .B(
        \b/SBOX[2].sbox/t[28] ), .Z(n1917) );
  XOR \b/SBOX[2].sbox/U107  ( .A(n1958), .B(n1918), .Z(n1963) );
  XOR \b/SBOX[2].sbox/U106  ( .A(\b/SBOX[2].sbox/t[5] ), .B(msg[20]), .Z(n1918) );
  XOR \b/SBOX[2].sbox/U105  ( .A(msg[23]), .B(n1919), .Z(n1959) );
  XOR \b/SBOX[2].sbox/U104  ( .A(\b/SBOX[2].sbox/t[7] ), .B(
        \b/SBOX[2].sbox/t[10] ), .Z(n1919) );
  XOR \b/SBOX[2].sbox/U103  ( .A(n1921), .B(n1920), .Z(\b/SBOX[2].sbox/t[42] )
         );
  XOR \b/SBOX[2].sbox/U102  ( .A(n1963), .B(n1959), .Z(n1920) );
  XOR \b/SBOX[2].sbox/U101  ( .A(\b/SBOX[2].sbox/t[28] ), .B(
        \b/SBOX[2].sbox/t[32] ), .Z(n1921) );
  XOR \b/SBOX[2].sbox/U100  ( .A(msg[17]), .B(n1922), .Z(n1961) );
  XOR \b/SBOX[2].sbox/U99  ( .A(msg[19]), .B(msg[18]), .Z(n1922) );
  XOR \b/SBOX[2].sbox/U98  ( .A(msg[21]), .B(n1961), .Z(\b/SBOX[2].sbox/y[16] ) );
  XOR \b/SBOX[2].sbox/U97  ( .A(\b/SBOX[2].sbox/y[16] ), .B(n1923), .Z(n1962)
         );
  XOR \b/SBOX[2].sbox/U96  ( .A(\b/SBOX[2].sbox/t[12] ), .B(
        \b/SBOX[2].sbox/t[15] ), .Z(n1923) );
  XOR \b/SBOX[2].sbox/U95  ( .A(n1962), .B(n1924), .Z(\b/SBOX[2].sbox/t[29] )
         );
  XOR \b/SBOX[2].sbox/U94  ( .A(\b/SBOX[2].sbox/t[28] ), .B(n1963), .Z(n1924)
         );
  XOR \b/SBOX[2].sbox/U93  ( .A(msg[16]), .B(n1925), .Z(\b/SBOX[2].sbox/y[1] )
         );
  XOR \b/SBOX[2].sbox/U92  ( .A(msg[22]), .B(msg[21]), .Z(n1925) );
  XOR \b/SBOX[2].sbox/U91  ( .A(msg[23]), .B(\b/SBOX[2].sbox/y[1] ), .Z(
        \b/SBOX[2].sbox/y[2] ) );
  XOR \b/SBOX[2].sbox/U90  ( .A(n1927), .B(n1926), .Z(\b/SBOX[2].sbox/t[25] )
         );
  XOR \b/SBOX[2].sbox/U89  ( .A(n1929), .B(n1928), .Z(n1926) );
  XOR \b/SBOX[2].sbox/U88  ( .A(msg[23]), .B(msg[21]), .Z(n1927) );
  XOR \b/SBOX[2].sbox/U87  ( .A(\b/SBOX[2].sbox/t[13] ), .B(
        \b/SBOX[2].sbox/t[15] ), .Z(n1928) );
  XOR \b/SBOX[2].sbox/U86  ( .A(\b/SBOX[2].sbox/t[3] ), .B(
        \b/SBOX[2].sbox/t[5] ), .Z(n1929) );
  XOR \b/SBOX[2].sbox/U85  ( .A(\b/SBOX[2].sbox/t[39] ), .B(
        \b/SBOX[2].sbox/t[25] ), .Z(\b/SBOX[2].sbox/t[40] ) );
  XOR \b/SBOX[2].sbox/U84  ( .A(msg[17]), .B(\b/SBOX[2].sbox/y[1] ), .Z(
        \b/SBOX[2].sbox/y[5] ) );
  XOR \b/SBOX[2].sbox/U83  ( .A(n1931), .B(n1930), .Z(\b/SBOX[2].sbox/y[15] )
         );
  XOR \b/SBOX[2].sbox/U82  ( .A(msg[19]), .B(msg[17]), .Z(n1930) );
  XOR \b/SBOX[2].sbox/U81  ( .A(msg[23]), .B(msg[20]), .Z(n1931) );
  XOR \b/SBOX[2].sbox/U80  ( .A(n1933), .B(n1932), .Z(\b/SBOX[2].sbox/t[21] )
         );
  XOR \b/SBOX[2].sbox/U79  ( .A(n1935), .B(n1934), .Z(n1932) );
  XOR \b/SBOX[2].sbox/U78  ( .A(\b/SBOX[2].sbox/y[15] ), .B(n1958), .Z(n1933)
         );
  XOR \b/SBOX[2].sbox/U77  ( .A(\b/SBOX[2].sbox/t[13] ), .B(msg[18]), .Z(n1934) );
  XOR \b/SBOX[2].sbox/U76  ( .A(\b/SBOX[2].sbox/t[3] ), .B(
        \b/SBOX[2].sbox/t[12] ), .Z(n1935) );
  XOR \b/SBOX[2].sbox/U75  ( .A(\b/SBOX[2].sbox/t[21] ), .B(n1936), .Z(
        \b/SBOX[2].sbox/t[43] ) );
  XOR \b/SBOX[2].sbox/U74  ( .A(\b/SBOX[2].sbox/t[28] ), .B(
        \b/SBOX[2].sbox/t[39] ), .Z(n1936) );
  XOR \b/SBOX[2].sbox/U73  ( .A(n1962), .B(n1959), .Z(\b/SBOX[2].sbox/t[24] )
         );
  XOR \b/SBOX[2].sbox/U72  ( .A(\b/SBOX[2].sbox/t[32] ), .B(
        \b/SBOX[2].sbox/t[24] ), .Z(\b/SBOX[2].sbox/t[33] ) );
  XOR \b/SBOX[2].sbox/U71  ( .A(msg[20]), .B(\b/SBOX[2].sbox/y[1] ), .Z(
        \b/SBOX[2].sbox/y[4] ) );
  XOR \b/SBOX[2].sbox/U70  ( .A(n1938), .B(n1937), .Z(\b/SBOX[2].sbox/t[30] )
         );
  XOR \b/SBOX[2].sbox/U69  ( .A(msg[17]), .B(n1939), .Z(n1937) );
  XOR \b/SBOX[2].sbox/U68  ( .A(\b/SBOX[2].sbox/t[13] ), .B(
        \b/SBOX[2].sbox/t[15] ), .Z(n1938) );
  XOR \b/SBOX[2].sbox/U67  ( .A(\b/SBOX[2].sbox/t[8] ), .B(
        \b/SBOX[2].sbox/t[10] ), .Z(n1939) );
  XOR \b/SBOX[2].sbox/U66  ( .A(\b/SBOX[2].sbox/t[30] ), .B(n1940), .Z(
        \b/SBOX[2].sbox/t[37] ) );
  XOR \b/SBOX[2].sbox/U65  ( .A(\b/SBOX[2].sbox/t[32] ), .B(
        \b/SBOX[2].sbox/t[36] ), .Z(n1940) );
  XOR \b/SBOX[2].sbox/U64  ( .A(msg[23]), .B(msg[18]), .Z(n1960) );
  XOR \b/SBOX[2].sbox/U63  ( .A(\b/SBOX[2].sbox/y[5] ), .B(n1960), .Z(
        \b/SBOX[2].sbox/y[3] ) );
  XOR \b/SBOX[2].sbox/U62  ( .A(n1942), .B(n1941), .Z(\b/SBOX[2].sbox/t[23] )
         );
  XOR \b/SBOX[2].sbox/U61  ( .A(n1944), .B(n1943), .Z(n1941) );
  XOR \b/SBOX[2].sbox/U60  ( .A(n1960), .B(n1945), .Z(n1942) );
  XOR \b/SBOX[2].sbox/U59  ( .A(msg[21]), .B(msg[19]), .Z(n1943) );
  XOR \b/SBOX[2].sbox/U58  ( .A(\b/SBOX[2].sbox/t[12] ), .B(
        \b/SBOX[2].sbox/t[13] ), .Z(n1944) );
  XOR \b/SBOX[2].sbox/U57  ( .A(\b/SBOX[2].sbox/t[7] ), .B(
        \b/SBOX[2].sbox/t[8] ), .Z(n1945) );
  XOR \b/SBOX[2].sbox/U56  ( .A(\b/SBOX[2].sbox/t[36] ), .B(
        \b/SBOX[2].sbox/t[23] ), .Z(\b/SBOX[2].sbox/t[44] ) );
  XOR \b/SBOX[2].sbox/U55  ( .A(n1960), .B(n1946), .Z(\b/SBOX[2].sbox/y[12] )
         );
  XOR \b/SBOX[2].sbox/U54  ( .A(msg[20]), .B(msg[17]), .Z(n1946) );
  XOR \b/SBOX[2].sbox/U53  ( .A(\b/SBOX[2].sbox/y[15] ), .B(n1947), .Z(
        \b/SBOX[2].sbox/y[10] ) );
  XOR \b/SBOX[2].sbox/U52  ( .A(msg[22]), .B(msg[21]), .Z(n1947) );
  XOR \b/SBOX[2].sbox/U51  ( .A(n1960), .B(n1948), .Z(\b/SBOX[2].sbox/y[17] )
         );
  XOR \b/SBOX[2].sbox/U50  ( .A(msg[21]), .B(msg[20]), .Z(n1948) );
  XOR \b/SBOX[2].sbox/U49  ( .A(msg[22]), .B(n1961), .Z(\b/SBOX[2].sbox/y[11] ) );
  XOR \b/SBOX[2].sbox/U48  ( .A(msg[16]), .B(\b/SBOX[2].sbox/y[11] ), .Z(
        \b/SBOX[2].sbox/y[7] ) );
  XOR \b/SBOX[2].sbox/U47  ( .A(msg[16]), .B(\b/SBOX[2].sbox/y[15] ), .Z(
        \b/SBOX[2].sbox/y[6] ) );
  XOR \b/SBOX[2].sbox/U46  ( .A(\b/SBOX[2].sbox/t[26] ), .B(
        \b/SBOX[2].sbox/t[24] ), .Z(\b/SBOX[2].sbox/t[27] ) );
  XOR \b/SBOX[2].sbox/U45  ( .A(\b/SBOX[2].sbox/t[36] ), .B(
        \b/SBOX[2].sbox/t[27] ), .Z(\b/SBOX[2].sbox/t[38] ) );
  XOR \b/SBOX[2].sbox/U44  ( .A(n1962), .B(n1949), .Z(\b/SBOX[2].sbox/t[31] )
         );
  XOR \b/SBOX[2].sbox/U43  ( .A(\b/SBOX[2].sbox/t[26] ), .B(n1963), .Z(n1949)
         );
  XOR \b/SBOX[1].sbox/U157  ( .A(\b/SBOX[1].sbox/z[12] ), .B(n1806), .Z(n1870)
         );
  XOR \b/SBOX[1].sbox/U156  ( .A(\b/SBOX[1].sbox/z[0] ), .B(
        \b/SBOX[1].sbox/z[2] ), .Z(n1806) );
  XOR \b/SBOX[1].sbox/U155  ( .A(n1808), .B(n1807), .Z(n1869) );
  XOR \b/SBOX[1].sbox/U154  ( .A(\b/SBOX[1].sbox/z[15] ), .B(
        \b/SBOX[1].sbox/z[16] ), .Z(n1807) );
  XOR \b/SBOX[1].sbox/U153  ( .A(\b/SBOX[1].sbox/z[5] ), .B(
        \b/SBOX[1].sbox/z[13] ), .Z(n1808) );
  XOR \b/SBOX[1].sbox/U152  ( .A(n1869), .B(n1809), .Z(n1883) );
  XOR \b/SBOX[1].sbox/U151  ( .A(\b/SBOX[1].sbox/z[3] ), .B(n1870), .Z(n1809)
         );
  XOR \b/SBOX[1].sbox/U150  ( .A(n1811), .B(n1810), .Z(n1884) );
  XOR \b/SBOX[1].sbox/U149  ( .A(n1869), .B(n1812), .Z(n1810) );
  XOR \b/SBOX[1].sbox/U148  ( .A(\b/SBOX[1].sbox/z[8] ), .B(
        \b/SBOX[1].sbox/z[12] ), .Z(n1811) );
  XOR \b/SBOX[1].sbox/U147  ( .A(\b/SBOX[1].sbox/z[4] ), .B(
        \b/SBOX[1].sbox/z[7] ), .Z(n1812) );
  XOR \b/SBOX[1].sbox/U146  ( .A(n1870), .B(n1813), .Z(n1872) );
  XOR \b/SBOX[1].sbox/U145  ( .A(\b/SBOX[1].sbox/z[8] ), .B(
        \b/SBOX[1].sbox/z[14] ), .Z(n1813) );
  XOR \b/SBOX[1].sbox/U144  ( .A(n1815), .B(n1814), .Z(n1885) );
  XOR \b/SBOX[1].sbox/U143  ( .A(\b/SBOX[1].sbox/z[17] ), .B(n1872), .Z(n1814)
         );
  XOR \b/SBOX[1].sbox/U142  ( .A(\b/SBOX[1].sbox/z[6] ), .B(
        \b/SBOX[1].sbox/z[15] ), .Z(n1815) );
  XOR \b/SBOX[1].sbox/U141  ( .A(\b/SBOX[1].sbox/z[9] ), .B(n1816), .Z(n1873)
         );
  XOR \b/SBOX[1].sbox/U140  ( .A(\b/SBOX[1].sbox/z[0] ), .B(
        \b/SBOX[1].sbox/z[1] ), .Z(n1816) );
  XOR \b/SBOX[1].sbox/U139  ( .A(\b/SBOX[1].sbox/z[16] ), .B(n1817), .Z(n1871)
         );
  XOR \b/SBOX[1].sbox/U138  ( .A(\b/SBOX[1].sbox/z[10] ), .B(
        \b/SBOX[1].sbox/z[15] ), .Z(n1817) );
  XOR \b/SBOX[1].sbox/U137  ( .A(n1819), .B(n1818), .Z(n1886) );
  XOR \b/SBOX[1].sbox/U136  ( .A(n1873), .B(n1871), .Z(n1818) );
  XOR \b/SBOX[1].sbox/U135  ( .A(\b/SBOX[1].sbox/z[6] ), .B(
        \b/SBOX[1].sbox/z[7] ), .Z(n1819) );
  XOR \b/SBOX[1].sbox/U134  ( .A(\b/SBOX[1].sbox/z[4] ), .B(n1871), .Z(n1874)
         );
  XOR \b/SBOX[1].sbox/U133  ( .A(n1874), .B(n1820), .Z(n1875) );
  XOR \b/SBOX[1].sbox/U132  ( .A(\b/SBOX[1].sbox/z[3] ), .B(
        \b/SBOX[1].sbox/z[7] ), .Z(n1820) );
  XOR \b/SBOX[1].sbox/U131  ( .A(n1872), .B(n1821), .Z(shift_row_out[106]) );
  XOR \b/SBOX[1].sbox/U130  ( .A(\b/SBOX[1].sbox/z[11] ), .B(n1875), .Z(n1821)
         );
  XOR \b/SBOX[1].sbox/U129  ( .A(n1823), .B(n1822), .Z(shift_row_out[107]) );
  XOR \b/SBOX[1].sbox/U128  ( .A(n1874), .B(n1824), .Z(n1822) );
  XOR \b/SBOX[1].sbox/U127  ( .A(\b/SBOX[1].sbox/z[5] ), .B(
        \b/SBOX[1].sbox/z[9] ), .Z(n1823) );
  XOR \b/SBOX[1].sbox/U126  ( .A(\b/SBOX[1].sbox/z[1] ), .B(
        \b/SBOX[1].sbox/z[2] ), .Z(n1824) );
  XOR \b/SBOX[1].sbox/U125  ( .A(n1873), .B(n1825), .Z(shift_row_out[108]) );
  XOR \b/SBOX[1].sbox/U124  ( .A(\b/SBOX[1].sbox/z[3] ), .B(n1874), .Z(n1825)
         );
  XOR \b/SBOX[1].sbox/U123  ( .A(n1875), .B(n1826), .Z(shift_row_out[111]) );
  XOR \b/SBOX[1].sbox/U122  ( .A(\b/SBOX[1].sbox/z[6] ), .B(
        \b/SBOX[1].sbox/z[9] ), .Z(n1826) );
  XOR \b/SBOX[1].sbox/U121  ( .A(n1828), .B(n1827), .Z(n1876) );
  XOR \b/SBOX[1].sbox/U120  ( .A(n1830), .B(n1829), .Z(n1827) );
  XOR \b/SBOX[1].sbox/U119  ( .A(msg[13]), .B(msg[9]), .Z(n1828) );
  XOR \b/SBOX[1].sbox/U118  ( .A(\b/SBOX[1].sbox/t[36] ), .B(
        \b/SBOX[1].sbox/t[39] ), .Z(n1829) );
  XOR \b/SBOX[1].sbox/U117  ( .A(\b/SBOX[1].sbox/t[3] ), .B(
        \b/SBOX[1].sbox/t[8] ), .Z(n1830) );
  XOR \b/SBOX[1].sbox/U116  ( .A(n1832), .B(n1831), .Z(\b/SBOX[1].sbox/t[41] )
         );
  XOR \b/SBOX[1].sbox/U115  ( .A(n1876), .B(n1833), .Z(n1831) );
  XOR \b/SBOX[1].sbox/U114  ( .A(\b/SBOX[1].sbox/t[32] ), .B(msg[15]), .Z(
        n1832) );
  XOR \b/SBOX[1].sbox/U113  ( .A(\b/SBOX[1].sbox/t[5] ), .B(
        \b/SBOX[1].sbox/t[10] ), .Z(n1833) );
  XOR \b/SBOX[1].sbox/U112  ( .A(\b/SBOX[1].sbox/t[2] ), .B(msg[14]), .Z(n1877) );
  XOR \b/SBOX[1].sbox/U111  ( .A(n1835), .B(n1834), .Z(\b/SBOX[1].sbox/t[45] )
         );
  XOR \b/SBOX[1].sbox/U110  ( .A(n1877), .B(n1836), .Z(n1834) );
  XOR \b/SBOX[1].sbox/U109  ( .A(msg[12]), .B(n1876), .Z(n1835) );
  XOR \b/SBOX[1].sbox/U108  ( .A(\b/SBOX[1].sbox/t[7] ), .B(
        \b/SBOX[1].sbox/t[28] ), .Z(n1836) );
  XOR \b/SBOX[1].sbox/U107  ( .A(n1877), .B(n1837), .Z(n1882) );
  XOR \b/SBOX[1].sbox/U106  ( .A(\b/SBOX[1].sbox/t[5] ), .B(msg[12]), .Z(n1837) );
  XOR \b/SBOX[1].sbox/U105  ( .A(msg[15]), .B(n1838), .Z(n1878) );
  XOR \b/SBOX[1].sbox/U104  ( .A(\b/SBOX[1].sbox/t[7] ), .B(
        \b/SBOX[1].sbox/t[10] ), .Z(n1838) );
  XOR \b/SBOX[1].sbox/U103  ( .A(n1840), .B(n1839), .Z(\b/SBOX[1].sbox/t[42] )
         );
  XOR \b/SBOX[1].sbox/U102  ( .A(n1882), .B(n1878), .Z(n1839) );
  XOR \b/SBOX[1].sbox/U101  ( .A(\b/SBOX[1].sbox/t[28] ), .B(
        \b/SBOX[1].sbox/t[32] ), .Z(n1840) );
  XOR \b/SBOX[1].sbox/U100  ( .A(msg[9]), .B(n1841), .Z(n1880) );
  XOR \b/SBOX[1].sbox/U99  ( .A(msg[11]), .B(msg[10]), .Z(n1841) );
  XOR \b/SBOX[1].sbox/U98  ( .A(msg[13]), .B(n1880), .Z(\b/SBOX[1].sbox/y[16] ) );
  XOR \b/SBOX[1].sbox/U97  ( .A(\b/SBOX[1].sbox/y[16] ), .B(n1842), .Z(n1881)
         );
  XOR \b/SBOX[1].sbox/U96  ( .A(\b/SBOX[1].sbox/t[12] ), .B(
        \b/SBOX[1].sbox/t[15] ), .Z(n1842) );
  XOR \b/SBOX[1].sbox/U95  ( .A(n1881), .B(n1843), .Z(\b/SBOX[1].sbox/t[29] )
         );
  XOR \b/SBOX[1].sbox/U94  ( .A(\b/SBOX[1].sbox/t[28] ), .B(n1882), .Z(n1843)
         );
  XOR \b/SBOX[1].sbox/U93  ( .A(msg[8]), .B(n1844), .Z(\b/SBOX[1].sbox/y[1] )
         );
  XOR \b/SBOX[1].sbox/U92  ( .A(msg[14]), .B(msg[13]), .Z(n1844) );
  XOR \b/SBOX[1].sbox/U91  ( .A(msg[15]), .B(\b/SBOX[1].sbox/y[1] ), .Z(
        \b/SBOX[1].sbox/y[2] ) );
  XOR \b/SBOX[1].sbox/U90  ( .A(n1846), .B(n1845), .Z(\b/SBOX[1].sbox/t[25] )
         );
  XOR \b/SBOX[1].sbox/U89  ( .A(n1848), .B(n1847), .Z(n1845) );
  XOR \b/SBOX[1].sbox/U88  ( .A(msg[15]), .B(msg[13]), .Z(n1846) );
  XOR \b/SBOX[1].sbox/U87  ( .A(\b/SBOX[1].sbox/t[13] ), .B(
        \b/SBOX[1].sbox/t[15] ), .Z(n1847) );
  XOR \b/SBOX[1].sbox/U86  ( .A(\b/SBOX[1].sbox/t[3] ), .B(
        \b/SBOX[1].sbox/t[5] ), .Z(n1848) );
  XOR \b/SBOX[1].sbox/U85  ( .A(\b/SBOX[1].sbox/t[39] ), .B(
        \b/SBOX[1].sbox/t[25] ), .Z(\b/SBOX[1].sbox/t[40] ) );
  XOR \b/SBOX[1].sbox/U84  ( .A(msg[9]), .B(\b/SBOX[1].sbox/y[1] ), .Z(
        \b/SBOX[1].sbox/y[5] ) );
  XOR \b/SBOX[1].sbox/U83  ( .A(n1850), .B(n1849), .Z(\b/SBOX[1].sbox/y[15] )
         );
  XOR \b/SBOX[1].sbox/U82  ( .A(msg[11]), .B(msg[9]), .Z(n1849) );
  XOR \b/SBOX[1].sbox/U81  ( .A(msg[15]), .B(msg[12]), .Z(n1850) );
  XOR \b/SBOX[1].sbox/U80  ( .A(n1852), .B(n1851), .Z(\b/SBOX[1].sbox/t[21] )
         );
  XOR \b/SBOX[1].sbox/U79  ( .A(n1854), .B(n1853), .Z(n1851) );
  XOR \b/SBOX[1].sbox/U78  ( .A(\b/SBOX[1].sbox/y[15] ), .B(n1877), .Z(n1852)
         );
  XOR \b/SBOX[1].sbox/U77  ( .A(\b/SBOX[1].sbox/t[13] ), .B(msg[10]), .Z(n1853) );
  XOR \b/SBOX[1].sbox/U76  ( .A(\b/SBOX[1].sbox/t[3] ), .B(
        \b/SBOX[1].sbox/t[12] ), .Z(n1854) );
  XOR \b/SBOX[1].sbox/U75  ( .A(\b/SBOX[1].sbox/t[21] ), .B(n1855), .Z(
        \b/SBOX[1].sbox/t[43] ) );
  XOR \b/SBOX[1].sbox/U74  ( .A(\b/SBOX[1].sbox/t[28] ), .B(
        \b/SBOX[1].sbox/t[39] ), .Z(n1855) );
  XOR \b/SBOX[1].sbox/U73  ( .A(n1881), .B(n1878), .Z(\b/SBOX[1].sbox/t[24] )
         );
  XOR \b/SBOX[1].sbox/U72  ( .A(\b/SBOX[1].sbox/t[32] ), .B(
        \b/SBOX[1].sbox/t[24] ), .Z(\b/SBOX[1].sbox/t[33] ) );
  XOR \b/SBOX[1].sbox/U71  ( .A(msg[12]), .B(\b/SBOX[1].sbox/y[1] ), .Z(
        \b/SBOX[1].sbox/y[4] ) );
  XOR \b/SBOX[1].sbox/U70  ( .A(n1857), .B(n1856), .Z(\b/SBOX[1].sbox/t[30] )
         );
  XOR \b/SBOX[1].sbox/U69  ( .A(msg[9]), .B(n1858), .Z(n1856) );
  XOR \b/SBOX[1].sbox/U68  ( .A(\b/SBOX[1].sbox/t[13] ), .B(
        \b/SBOX[1].sbox/t[15] ), .Z(n1857) );
  XOR \b/SBOX[1].sbox/U67  ( .A(\b/SBOX[1].sbox/t[8] ), .B(
        \b/SBOX[1].sbox/t[10] ), .Z(n1858) );
  XOR \b/SBOX[1].sbox/U66  ( .A(\b/SBOX[1].sbox/t[30] ), .B(n1859), .Z(
        \b/SBOX[1].sbox/t[37] ) );
  XOR \b/SBOX[1].sbox/U65  ( .A(\b/SBOX[1].sbox/t[32] ), .B(
        \b/SBOX[1].sbox/t[36] ), .Z(n1859) );
  XOR \b/SBOX[1].sbox/U64  ( .A(msg[15]), .B(msg[10]), .Z(n1879) );
  XOR \b/SBOX[1].sbox/U63  ( .A(\b/SBOX[1].sbox/y[5] ), .B(n1879), .Z(
        \b/SBOX[1].sbox/y[3] ) );
  XOR \b/SBOX[1].sbox/U62  ( .A(n1861), .B(n1860), .Z(\b/SBOX[1].sbox/t[23] )
         );
  XOR \b/SBOX[1].sbox/U61  ( .A(n1863), .B(n1862), .Z(n1860) );
  XOR \b/SBOX[1].sbox/U60  ( .A(n1879), .B(n1864), .Z(n1861) );
  XOR \b/SBOX[1].sbox/U59  ( .A(msg[13]), .B(msg[11]), .Z(n1862) );
  XOR \b/SBOX[1].sbox/U58  ( .A(\b/SBOX[1].sbox/t[12] ), .B(
        \b/SBOX[1].sbox/t[13] ), .Z(n1863) );
  XOR \b/SBOX[1].sbox/U57  ( .A(\b/SBOX[1].sbox/t[7] ), .B(
        \b/SBOX[1].sbox/t[8] ), .Z(n1864) );
  XOR \b/SBOX[1].sbox/U56  ( .A(\b/SBOX[1].sbox/t[36] ), .B(
        \b/SBOX[1].sbox/t[23] ), .Z(\b/SBOX[1].sbox/t[44] ) );
  XOR \b/SBOX[1].sbox/U55  ( .A(n1879), .B(n1865), .Z(\b/SBOX[1].sbox/y[12] )
         );
  XOR \b/SBOX[1].sbox/U54  ( .A(msg[12]), .B(msg[9]), .Z(n1865) );
  XOR \b/SBOX[1].sbox/U53  ( .A(\b/SBOX[1].sbox/y[15] ), .B(n1866), .Z(
        \b/SBOX[1].sbox/y[10] ) );
  XOR \b/SBOX[1].sbox/U52  ( .A(msg[14]), .B(msg[13]), .Z(n1866) );
  XOR \b/SBOX[1].sbox/U51  ( .A(n1879), .B(n1867), .Z(\b/SBOX[1].sbox/y[17] )
         );
  XOR \b/SBOX[1].sbox/U50  ( .A(msg[13]), .B(msg[12]), .Z(n1867) );
  XOR \b/SBOX[1].sbox/U49  ( .A(msg[14]), .B(n1880), .Z(\b/SBOX[1].sbox/y[11] ) );
  XOR \b/SBOX[1].sbox/U48  ( .A(msg[8]), .B(\b/SBOX[1].sbox/y[11] ), .Z(
        \b/SBOX[1].sbox/y[7] ) );
  XOR \b/SBOX[1].sbox/U47  ( .A(msg[8]), .B(\b/SBOX[1].sbox/y[15] ), .Z(
        \b/SBOX[1].sbox/y[6] ) );
  XOR \b/SBOX[1].sbox/U46  ( .A(\b/SBOX[1].sbox/t[26] ), .B(
        \b/SBOX[1].sbox/t[24] ), .Z(\b/SBOX[1].sbox/t[27] ) );
  XOR \b/SBOX[1].sbox/U45  ( .A(\b/SBOX[1].sbox/t[36] ), .B(
        \b/SBOX[1].sbox/t[27] ), .Z(\b/SBOX[1].sbox/t[38] ) );
  XOR \b/SBOX[1].sbox/U44  ( .A(n1881), .B(n1868), .Z(\b/SBOX[1].sbox/t[31] )
         );
  XOR \b/SBOX[1].sbox/U43  ( .A(\b/SBOX[1].sbox/t[26] ), .B(n1882), .Z(n1868)
         );
  XNOR U659 ( .A(n2939), .B(n2048), .Z(n1012) );
  XOR U660 ( .A(n2938), .B(n2047), .Z(n1021) );
  XOR U661 ( .A(\e/w[3][2] ), .B(nextKey[66]), .Z(n550) );
  MUX U662 ( .IN0(counter[0]), .IN1(n528), .SEL(counter[3]), .F(n1696) );
  IV U663 ( .A(counter[1]), .Z(n528) );
  XNOR U664 ( .A(n2694), .B(n2775), .Z(n1476) );
  XOR U665 ( .A(n2693), .B(n2774), .Z(n1485) );
  XNOR U666 ( .A(n2696), .B(n2291), .Z(n1513) );
  XOR U667 ( .A(n2937), .B(n2046), .Z(n1061) );
  XOR U668 ( .A(n2936), .B(n2045), .Z(n1082) );
  XNOR U669 ( .A(\b/SBOX[0].sbox/n91 ), .B(n3020), .Z(n1238) );
  XOR U670 ( .A(n1885), .B(n2776), .Z(n1531) );
  XNOR U671 ( .A(n1106), .B(n1012), .Z(n1105) );
  XNOR U672 ( .A(n564), .B(n563), .Z(n562) );
  XNOR U673 ( .A(\e/w[3][31] ), .B(\e/n291 ), .Z(nextKey[127]) );
  XNOR U674 ( .A(\e/w[3][30] ), .B(\e/n290 ), .Z(nextKey[126]) );
  XNOR U675 ( .A(\e/w[3][29] ), .B(\e/n289 ), .Z(nextKey[125]) );
  XNOR U676 ( .A(\e/w[3][28] ), .B(\e/n288 ), .Z(nextKey[124]) );
  XNOR U677 ( .A(\e/w[3][27] ), .B(\e/n287 ), .Z(nextKey[123]) );
  XNOR U678 ( .A(\e/w[3][26] ), .B(\e/n286 ), .Z(nextKey[122]) );
  XNOR U679 ( .A(\e/w[3][25] ), .B(\e/n285 ), .Z(nextKey[121]) );
  XNOR U680 ( .A(\e/w[3][23] ), .B(\e/n283 ), .Z(nextKey[119]) );
  XNOR U681 ( .A(\e/w[3][22] ), .B(\e/n282 ), .Z(nextKey[118]) );
  XNOR U682 ( .A(\e/w[3][21] ), .B(\e/n281 ), .Z(nextKey[117]) );
  XNOR U683 ( .A(\e/w[3][20] ), .B(\e/n280 ), .Z(nextKey[116]) );
  XNOR U684 ( .A(\e/w[3][19] ), .B(\e/n279 ), .Z(nextKey[115]) );
  XNOR U685 ( .A(\e/w[3][18] ), .B(\e/n278 ), .Z(nextKey[114]) );
  XNOR U686 ( .A(\e/w[3][17] ), .B(\e/n277 ), .Z(nextKey[113]) );
  XNOR U687 ( .A(\e/w[3][15] ), .B(\e/n275 ), .Z(nextKey[111]) );
  XNOR U688 ( .A(\e/w[3][14] ), .B(\e/n274 ), .Z(nextKey[110]) );
  XNOR U689 ( .A(\e/w[3][13] ), .B(\e/n273 ), .Z(nextKey[109]) );
  XNOR U690 ( .A(\e/w[3][12] ), .B(\e/n272 ), .Z(nextKey[108]) );
  XNOR U691 ( .A(\e/w[3][11] ), .B(\e/n271 ), .Z(nextKey[107]) );
  XNOR U692 ( .A(\e/w[3][10] ), .B(\e/n270 ), .Z(nextKey[106]) );
  XNOR U693 ( .A(\e/w[3][9] ), .B(\e/n269 ), .Z(nextKey[105]) );
  XOR U694 ( .A(\e/w[3][7] ), .B(nextKey[71]), .Z(n545) );
  XOR U695 ( .A(\e/w[3][6] ), .B(nextKey[70]), .Z(n546) );
  XOR U696 ( .A(\e/w[3][5] ), .B(nextKey[69]), .Z(n547) );
  XOR U697 ( .A(\e/w[3][4] ), .B(nextKey[68]), .Z(n548) );
  XOR U698 ( .A(\e/w[3][3] ), .B(nextKey[67]), .Z(n549) );
  XOR U699 ( .A(\e/w[3][1] ), .B(nextKey[65]), .Z(n551) );
  MUX U700 ( .IN0(n1703), .IN1(counter[3]), .SEL(counter[0]), .F(n1701) );
  XNOR U701 ( .A(n3265), .B(n3264), .Z(n529) );
  XNOR U702 ( .A(n3261), .B(n3260), .Z(n530) );
  XNOR U703 ( .A(n3257), .B(n3256), .Z(n531) );
  XNOR U704 ( .A(n3315), .B(n3255), .Z(n532) );
  XNOR U705 ( .A(n3188), .B(n3187), .Z(n533) );
  XNOR U706 ( .A(n3184), .B(n3183), .Z(n534) );
  XNOR U707 ( .A(n3180), .B(n3179), .Z(n535) );
  XNOR U708 ( .A(n3238), .B(n3178), .Z(n536) );
  XNOR U709 ( .A(n3111), .B(n3110), .Z(n537) );
  XNOR U710 ( .A(n3107), .B(n3106), .Z(n538) );
  XNOR U711 ( .A(n3103), .B(n3102), .Z(n539) );
  XNOR U712 ( .A(n3161), .B(n3101), .Z(n540) );
  XNOR U713 ( .A(n3034), .B(n3033), .Z(n541) );
  XNOR U714 ( .A(n3030), .B(n3029), .Z(n542) );
  XNOR U715 ( .A(n3026), .B(n3025), .Z(n543) );
  XNOR U716 ( .A(n3084), .B(n3024), .Z(n544) );
  XNOR U717 ( .A(\e/n74 ), .B(nextKey[64]), .Z(n552) );
  XOR U718 ( .A(n553), .B(key[9]), .Z(o[9]) );
  NAND U719 ( .A(n554), .B(n555), .Z(n553) );
  NAND U720 ( .A(n556), .B(msg[9]), .Z(n555) );
  AND U721 ( .A(n557), .B(n558), .Z(n554) );
  NAND U722 ( .A(n559), .B(n560), .Z(n558) );
  XOR U723 ( .A(n561), .B(n562), .Z(n559) );
  XOR U724 ( .A(n2613), .B(n565), .Z(n561) );
  NANDN U725 ( .B(n2208), .A(n566), .Z(n557) );
  XOR U726 ( .A(n567), .B(key[99]), .Z(o[99]) );
  NAND U727 ( .A(n568), .B(n569), .Z(n567) );
  NAND U728 ( .A(n556), .B(msg[99]), .Z(n569) );
  AND U729 ( .A(n570), .B(n571), .Z(n568) );
  NAND U730 ( .A(n572), .B(n560), .Z(n571) );
  XOR U731 ( .A(n573), .B(n574), .Z(n572) );
  XOR U732 ( .A(n575), .B(n576), .Z(n574) );
  XOR U733 ( .A(shift_row_out[106]), .B(n577), .Z(n573) );
  XOR U734 ( .A(shift_row_out[98]), .B(shift_row_out[107]), .Z(n577) );
  NAND U735 ( .A(n566), .B(shift_row_out[99]), .Z(n570) );
  XOR U736 ( .A(n578), .B(key[98]), .Z(o[98]) );
  NAND U737 ( .A(n579), .B(n580), .Z(n578) );
  NAND U738 ( .A(n556), .B(msg[98]), .Z(n580) );
  AND U739 ( .A(n581), .B(n582), .Z(n579) );
  NAND U740 ( .A(n583), .B(n560), .Z(n582) );
  XOR U741 ( .A(n584), .B(n585), .Z(n583) );
  XNOR U742 ( .A(n2775), .B(n586), .Z(n585) );
  XNOR U743 ( .A(shift_row_out[106]), .B(n587), .Z(n584) );
  NAND U744 ( .A(n566), .B(shift_row_out[98]), .Z(n581) );
  XOR U745 ( .A(n588), .B(key[97]), .Z(o[97]) );
  NAND U746 ( .A(n589), .B(n590), .Z(n588) );
  NAND U747 ( .A(n556), .B(msg[97]), .Z(n590) );
  AND U748 ( .A(n591), .B(n592), .Z(n589) );
  NAND U749 ( .A(n593), .B(n560), .Z(n592) );
  XOR U750 ( .A(n594), .B(n595), .Z(n593) );
  XOR U751 ( .A(n575), .B(n596), .Z(n595) );
  XNOR U752 ( .A(n2774), .B(n597), .Z(n594) );
  XNOR U753 ( .A(n587), .B(n1883), .Z(n597) );
  NANDN U754 ( .B(n2775), .A(n566), .Z(n591) );
  XOR U755 ( .A(n598), .B(key[96]), .Z(o[96]) );
  NAND U756 ( .A(n599), .B(n600), .Z(n598) );
  NAND U757 ( .A(n556), .B(msg[96]), .Z(n600) );
  AND U758 ( .A(n601), .B(n602), .Z(n599) );
  NAND U759 ( .A(n603), .B(n560), .Z(n602) );
  XNOR U760 ( .A(n604), .B(n605), .Z(n603) );
  XOR U761 ( .A(n1883), .B(n575), .Z(n604) );
  IV U762 ( .A(n606), .Z(n575) );
  NANDN U763 ( .B(n2774), .A(n566), .Z(n601) );
  XOR U764 ( .A(n607), .B(key[95]), .Z(o[95]) );
  NAND U765 ( .A(n608), .B(n609), .Z(n607) );
  NAND U766 ( .A(n556), .B(msg[95]), .Z(n609) );
  AND U767 ( .A(n610), .B(n611), .Z(n608) );
  NAND U768 ( .A(n612), .B(n560), .Z(n611) );
  XOR U769 ( .A(n613), .B(n614), .Z(n612) );
  XNOR U770 ( .A(n2372), .B(n615), .Z(n614) );
  XOR U771 ( .A(shift_row_out[71]), .B(n2453), .Z(n613) );
  NAND U772 ( .A(n566), .B(shift_row_out[95]), .Z(n610) );
  XOR U773 ( .A(n616), .B(key[94]), .Z(o[94]) );
  NAND U774 ( .A(n617), .B(n618), .Z(n616) );
  NAND U775 ( .A(n556), .B(msg[94]), .Z(n618) );
  AND U776 ( .A(n619), .B(n620), .Z(n617) );
  NAND U777 ( .A(n621), .B(n560), .Z(n620) );
  XOR U778 ( .A(n622), .B(n623), .Z(n621) );
  XNOR U779 ( .A(n2453), .B(n624), .Z(n623) );
  XOR U780 ( .A(n2371), .B(n625), .Z(n622) );
  NANDN U781 ( .B(n2372), .A(n566), .Z(n619) );
  XOR U782 ( .A(n626), .B(key[93]), .Z(o[93]) );
  NAND U783 ( .A(n627), .B(n628), .Z(n626) );
  NAND U784 ( .A(n556), .B(msg[93]), .Z(n628) );
  AND U785 ( .A(n629), .B(n630), .Z(n627) );
  NAND U786 ( .A(n631), .B(n560), .Z(n630) );
  XOR U787 ( .A(n632), .B(n633), .Z(n631) );
  XOR U788 ( .A(shift_row_out[92]), .B(shift_row_out[68]), .Z(n633) );
  XOR U789 ( .A(n2452), .B(n634), .Z(n632) );
  NANDN U790 ( .B(n2371), .A(n566), .Z(n629) );
  XOR U791 ( .A(n635), .B(key[92]), .Z(o[92]) );
  NAND U792 ( .A(n636), .B(n637), .Z(n635) );
  NAND U793 ( .A(n556), .B(msg[92]), .Z(n637) );
  AND U794 ( .A(n638), .B(n639), .Z(n636) );
  NAND U795 ( .A(n640), .B(n560), .Z(n639) );
  XOR U796 ( .A(n641), .B(n642), .Z(n640) );
  XOR U797 ( .A(n643), .B(n644), .Z(n642) );
  XOR U798 ( .A(shift_row_out[67]), .B(n645), .Z(n641) );
  XOR U799 ( .A(shift_row_out[91]), .B(shift_row_out[68]), .Z(n645) );
  NAND U800 ( .A(n566), .B(shift_row_out[92]), .Z(n638) );
  XOR U801 ( .A(n646), .B(key[91]), .Z(o[91]) );
  NAND U802 ( .A(n647), .B(n648), .Z(n646) );
  NAND U803 ( .A(n556), .B(msg[91]), .Z(n648) );
  AND U804 ( .A(n649), .B(n650), .Z(n647) );
  NAND U805 ( .A(n651), .B(n560), .Z(n650) );
  XOR U806 ( .A(n652), .B(n653), .Z(n651) );
  XOR U807 ( .A(n643), .B(n654), .Z(n653) );
  XOR U808 ( .A(shift_row_out[66]), .B(n655), .Z(n652) );
  XOR U809 ( .A(shift_row_out[90]), .B(shift_row_out[67]), .Z(n655) );
  NAND U810 ( .A(n566), .B(shift_row_out[91]), .Z(n649) );
  XOR U811 ( .A(n656), .B(key[90]), .Z(o[90]) );
  NAND U812 ( .A(n657), .B(n658), .Z(n656) );
  NAND U813 ( .A(msg[90]), .B(n556), .Z(n658) );
  AND U814 ( .A(n659), .B(n660), .Z(n657) );
  NAND U815 ( .A(n661), .B(n560), .Z(n660) );
  XOR U816 ( .A(n662), .B(n663), .Z(n661) );
  XNOR U817 ( .A(n2370), .B(n664), .Z(n663) );
  XOR U818 ( .A(shift_row_out[66]), .B(n2451), .Z(n662) );
  NAND U819 ( .A(n566), .B(shift_row_out[90]), .Z(n659) );
  XOR U820 ( .A(n665), .B(key[8]), .Z(o[8]) );
  NAND U821 ( .A(n666), .B(n667), .Z(n665) );
  NAND U822 ( .A(n556), .B(msg[8]), .Z(n667) );
  AND U823 ( .A(n668), .B(n669), .Z(n666) );
  NAND U824 ( .A(n670), .B(n560), .Z(n669) );
  XNOR U825 ( .A(n671), .B(n672), .Z(n670) );
  XNOR U826 ( .A(\b/SBOX[0].sbox/n88 ), .B(n564), .Z(n671) );
  NANDN U827 ( .B(n2207), .A(n566), .Z(n668) );
  XOR U828 ( .A(n673), .B(key[89]), .Z(o[89]) );
  NAND U829 ( .A(n674), .B(n675), .Z(n673) );
  NAND U830 ( .A(n556), .B(msg[89]), .Z(n675) );
  AND U831 ( .A(n676), .B(n677), .Z(n674) );
  NAND U832 ( .A(n678), .B(n560), .Z(n677) );
  XOR U833 ( .A(n679), .B(n680), .Z(n678) );
  XOR U834 ( .A(n643), .B(n681), .Z(n680) );
  XNOR U835 ( .A(n2369), .B(n682), .Z(n679) );
  XNOR U836 ( .A(n2451), .B(n683), .Z(n682) );
  NANDN U837 ( .B(n2370), .A(n566), .Z(n676) );
  XOR U838 ( .A(n684), .B(key[88]), .Z(o[88]) );
  NAND U839 ( .A(n685), .B(n686), .Z(n684) );
  NAND U840 ( .A(n556), .B(msg[88]), .Z(n686) );
  AND U841 ( .A(n687), .B(n688), .Z(n685) );
  NAND U842 ( .A(n689), .B(n560), .Z(n688) );
  XNOR U843 ( .A(n690), .B(n691), .Z(n689) );
  XOR U844 ( .A(n2450), .B(n643), .Z(n690) );
  XNOR U845 ( .A(shift_row_out[71]), .B(shift_row_out[95]), .Z(n643) );
  NANDN U846 ( .B(n2369), .A(n566), .Z(n687) );
  XOR U847 ( .A(n692), .B(key[87]), .Z(o[87]) );
  NAND U848 ( .A(n693), .B(n694), .Z(n692) );
  NAND U849 ( .A(n556), .B(msg[87]), .Z(n694) );
  AND U850 ( .A(n695), .B(n696), .Z(n693) );
  NAND U851 ( .A(n697), .B(n560), .Z(n696) );
  XOR U852 ( .A(n698), .B(n699), .Z(n697) );
  XNOR U853 ( .A(shift_row_out[71]), .B(n700), .Z(n699) );
  XNOR U854 ( .A(shift_row_out[95]), .B(n701), .Z(n698) );
  NAND U855 ( .A(n566), .B(shift_row_out[87]), .Z(n695) );
  XOR U856 ( .A(n702), .B(key[86]), .Z(o[86]) );
  NAND U857 ( .A(n703), .B(n704), .Z(n702) );
  NAND U858 ( .A(n556), .B(msg[86]), .Z(n704) );
  AND U859 ( .A(n705), .B(n706), .Z(n703) );
  NAND U860 ( .A(n707), .B(n560), .Z(n706) );
  XOR U861 ( .A(n708), .B(n709), .Z(n707) );
  XOR U862 ( .A(n2453), .B(n2372), .Z(n709) );
  XNOR U863 ( .A(n710), .B(n711), .Z(n708) );
  NANDN U864 ( .B(n1967), .A(n566), .Z(n705) );
  XOR U865 ( .A(n712), .B(key[85]), .Z(o[85]) );
  NAND U866 ( .A(n713), .B(n714), .Z(n712) );
  NAND U867 ( .A(n556), .B(msg[85]), .Z(n714) );
  AND U868 ( .A(n715), .B(n716), .Z(n713) );
  NAND U869 ( .A(n717), .B(n560), .Z(n716) );
  XOR U870 ( .A(n718), .B(n719), .Z(n717) );
  XNOR U871 ( .A(n624), .B(n2371), .Z(n719) );
  XNOR U872 ( .A(n720), .B(n721), .Z(n718) );
  NANDN U873 ( .B(n1966), .A(n566), .Z(n715) );
  XOR U874 ( .A(n722), .B(key[84]), .Z(o[84]) );
  NAND U875 ( .A(n723), .B(n724), .Z(n722) );
  NAND U876 ( .A(n556), .B(msg[84]), .Z(n724) );
  AND U877 ( .A(n725), .B(n726), .Z(n723) );
  NAND U878 ( .A(n727), .B(n560), .Z(n726) );
  XOR U879 ( .A(n728), .B(n729), .Z(n727) );
  XOR U880 ( .A(n730), .B(n731), .Z(n729) );
  XOR U881 ( .A(shift_row_out[68]), .B(n732), .Z(n728) );
  XOR U882 ( .A(shift_row_out[92]), .B(shift_row_out[76]), .Z(n732) );
  NAND U883 ( .A(n566), .B(shift_row_out[84]), .Z(n725) );
  XOR U884 ( .A(n733), .B(key[83]), .Z(o[83]) );
  NAND U885 ( .A(n734), .B(n735), .Z(n733) );
  NAND U886 ( .A(n556), .B(msg[83]), .Z(n735) );
  AND U887 ( .A(n736), .B(n737), .Z(n734) );
  NAND U888 ( .A(n738), .B(n560), .Z(n737) );
  XOR U889 ( .A(n739), .B(n740), .Z(n738) );
  XOR U890 ( .A(n731), .B(n741), .Z(n740) );
  XOR U891 ( .A(shift_row_out[67]), .B(n742), .Z(n739) );
  XOR U892 ( .A(shift_row_out[91]), .B(shift_row_out[75]), .Z(n742) );
  NAND U893 ( .A(n566), .B(shift_row_out[83]), .Z(n736) );
  XOR U894 ( .A(n743), .B(key[82]), .Z(o[82]) );
  NAND U895 ( .A(n744), .B(n745), .Z(n743) );
  NAND U896 ( .A(msg[82]), .B(n556), .Z(n745) );
  AND U897 ( .A(n746), .B(n747), .Z(n744) );
  NAND U898 ( .A(n748), .B(n560), .Z(n747) );
  XOR U899 ( .A(n749), .B(n750), .Z(n748) );
  XNOR U900 ( .A(shift_row_out[66]), .B(n751), .Z(n750) );
  XOR U901 ( .A(shift_row_out[90]), .B(shift_row_out[74]), .Z(n749) );
  NAND U902 ( .A(n566), .B(shift_row_out[82]), .Z(n746) );
  XOR U903 ( .A(n752), .B(key[81]), .Z(o[81]) );
  NAND U904 ( .A(n753), .B(n754), .Z(n752) );
  NAND U905 ( .A(n556), .B(msg[81]), .Z(n754) );
  AND U906 ( .A(n755), .B(n756), .Z(n753) );
  NAND U907 ( .A(n757), .B(n560), .Z(n756) );
  XOR U908 ( .A(n758), .B(n759), .Z(n757) );
  XOR U909 ( .A(n731), .B(n760), .Z(n759) );
  XNOR U910 ( .A(n2856), .B(n761), .Z(n758) );
  XOR U911 ( .A(n2451), .B(n2370), .Z(n761) );
  NANDN U912 ( .B(n1965), .A(n566), .Z(n755) );
  XOR U913 ( .A(n762), .B(key[80]), .Z(o[80]) );
  NAND U914 ( .A(n763), .B(n764), .Z(n762) );
  NAND U915 ( .A(n556), .B(msg[80]), .Z(n764) );
  AND U916 ( .A(n765), .B(n766), .Z(n763) );
  NAND U917 ( .A(n767), .B(n560), .Z(n766) );
  XOR U918 ( .A(n768), .B(n769), .Z(n767) );
  XNOR U919 ( .A(n683), .B(n2369), .Z(n769) );
  XOR U920 ( .A(n2855), .B(n731), .Z(n768) );
  NANDN U921 ( .B(n1964), .A(n566), .Z(n765) );
  XOR U922 ( .A(n770), .B(key[7]), .Z(o[7]) );
  NAND U923 ( .A(n771), .B(n772), .Z(n770) );
  NAND U924 ( .A(n556), .B(msg[7]), .Z(n772) );
  AND U925 ( .A(n773), .B(n774), .Z(n771) );
  NAND U926 ( .A(n775), .B(n560), .Z(n774) );
  XOR U927 ( .A(n776), .B(n777), .Z(n775) );
  XOR U928 ( .A(\b/SBOX[0].sbox/n91 ), .B(n778), .Z(n777) );
  XNOR U929 ( .A(shift_row_out[15]), .B(n779), .Z(n776) );
  NAND U930 ( .A(n566), .B(shift_row_out[7]), .Z(n773) );
  XOR U931 ( .A(n780), .B(key[79]), .Z(o[79]) );
  NAND U932 ( .A(n781), .B(n782), .Z(n780) );
  NAND U933 ( .A(n556), .B(msg[79]), .Z(n782) );
  AND U934 ( .A(n783), .B(n784), .Z(n781) );
  NAND U935 ( .A(n785), .B(n560), .Z(n784) );
  XNOR U936 ( .A(n731), .B(n786), .Z(n785) );
  XNOR U937 ( .A(shift_row_out[71]), .B(n625), .Z(n786) );
  XOR U938 ( .A(n2858), .B(n787), .Z(n625) );
  NANDN U939 ( .B(n701), .A(n566), .Z(n783) );
  XOR U940 ( .A(n788), .B(key[78]), .Z(o[78]) );
  NAND U941 ( .A(n789), .B(n790), .Z(n788) );
  NAND U942 ( .A(n556), .B(msg[78]), .Z(n790) );
  AND U943 ( .A(n791), .B(n792), .Z(n789) );
  NAND U944 ( .A(n793), .B(n560), .Z(n792) );
  XNOR U945 ( .A(n794), .B(n700), .Z(n793) );
  XOR U946 ( .A(n2453), .B(n634), .Z(n794) );
  XOR U947 ( .A(n2857), .B(n795), .Z(n634) );
  NANDN U948 ( .B(n2858), .A(n566), .Z(n791) );
  XOR U949 ( .A(n796), .B(key[77]), .Z(o[77]) );
  NAND U950 ( .A(n797), .B(n798), .Z(n796) );
  NAND U951 ( .A(n556), .B(msg[77]), .Z(n798) );
  AND U952 ( .A(n799), .B(n800), .Z(n797) );
  NAND U953 ( .A(n801), .B(n560), .Z(n800) );
  XNOR U954 ( .A(n802), .B(n711), .Z(n801) );
  XOR U955 ( .A(n2452), .B(n644), .Z(n802) );
  XNOR U956 ( .A(shift_row_out[76]), .B(shift_row_out[84]), .Z(n644) );
  NANDN U957 ( .B(n2857), .A(n566), .Z(n799) );
  XOR U958 ( .A(n803), .B(key[76]), .Z(o[76]) );
  NAND U959 ( .A(n804), .B(n805), .Z(n803) );
  NAND U960 ( .A(n556), .B(msg[76]), .Z(n805) );
  AND U961 ( .A(n806), .B(n807), .Z(n804) );
  NAND U962 ( .A(n808), .B(n560), .Z(n807) );
  XOR U963 ( .A(n809), .B(n810), .Z(n808) );
  XOR U964 ( .A(n654), .B(n721), .Z(n810) );
  XNOR U965 ( .A(shift_row_out[75]), .B(shift_row_out[83]), .Z(n654) );
  XNOR U966 ( .A(shift_row_out[68]), .B(n615), .Z(n809) );
  NAND U967 ( .A(n566), .B(shift_row_out[76]), .Z(n806) );
  XOR U968 ( .A(n811), .B(key[75]), .Z(o[75]) );
  NAND U969 ( .A(n812), .B(n813), .Z(n811) );
  NAND U970 ( .A(n556), .B(msg[75]), .Z(n813) );
  AND U971 ( .A(n814), .B(n815), .Z(n812) );
  NAND U972 ( .A(n816), .B(n560), .Z(n815) );
  XOR U973 ( .A(n817), .B(n818), .Z(n816) );
  XOR U974 ( .A(n664), .B(n730), .Z(n818) );
  XNOR U975 ( .A(shift_row_out[74]), .B(shift_row_out[82]), .Z(n664) );
  XNOR U976 ( .A(shift_row_out[67]), .B(n615), .Z(n817) );
  NAND U977 ( .A(n566), .B(shift_row_out[75]), .Z(n814) );
  XOR U978 ( .A(n819), .B(key[74]), .Z(o[74]) );
  NAND U979 ( .A(n820), .B(n821), .Z(n819) );
  NAND U980 ( .A(msg[74]), .B(n556), .Z(n821) );
  AND U981 ( .A(n822), .B(n823), .Z(n820) );
  NAND U982 ( .A(n824), .B(n560), .Z(n823) );
  XNOR U983 ( .A(n741), .B(n825), .Z(n824) );
  XNOR U984 ( .A(shift_row_out[66]), .B(n681), .Z(n825) );
  XNOR U985 ( .A(n2856), .B(n1965), .Z(n681) );
  NAND U986 ( .A(n566), .B(shift_row_out[74]), .Z(n822) );
  XOR U987 ( .A(n826), .B(key[73]), .Z(o[73]) );
  NAND U988 ( .A(n827), .B(n828), .Z(n826) );
  NAND U989 ( .A(n556), .B(msg[73]), .Z(n828) );
  AND U990 ( .A(n829), .B(n830), .Z(n827) );
  NAND U991 ( .A(n831), .B(n560), .Z(n830) );
  XOR U992 ( .A(n832), .B(n833), .Z(n831) );
  XOR U993 ( .A(n691), .B(n751), .Z(n833) );
  XNOR U994 ( .A(n2855), .B(n1964), .Z(n691) );
  XOR U995 ( .A(n2451), .B(n615), .Z(n832) );
  NANDN U996 ( .B(n2856), .A(n566), .Z(n829) );
  XOR U997 ( .A(n834), .B(key[72]), .Z(o[72]) );
  NAND U998 ( .A(n835), .B(n836), .Z(n834) );
  NAND U999 ( .A(n556), .B(msg[72]), .Z(n836) );
  AND U1000 ( .A(n837), .B(n838), .Z(n835) );
  NAND U1001 ( .A(n839), .B(n560), .Z(n838) );
  XNOR U1002 ( .A(n840), .B(n760), .Z(n839) );
  XOR U1003 ( .A(n2450), .B(n615), .Z(n840) );
  XNOR U1004 ( .A(shift_row_out[79]), .B(shift_row_out[87]), .Z(n615) );
  NANDN U1005 ( .B(n2855), .A(n566), .Z(n837) );
  XOR U1006 ( .A(n841), .B(key[71]), .Z(o[71]) );
  NAND U1007 ( .A(n842), .B(n843), .Z(n841) );
  NAND U1008 ( .A(n556), .B(msg[71]), .Z(n843) );
  AND U1009 ( .A(n844), .B(n845), .Z(n842) );
  NAND U1010 ( .A(n846), .B(n560), .Z(n845) );
  XOR U1011 ( .A(n847), .B(n848), .Z(n846) );
  XOR U1012 ( .A(n710), .B(n731), .Z(n848) );
  XNOR U1013 ( .A(shift_row_out[87]), .B(shift_row_out[95]), .Z(n731) );
  IV U1014 ( .A(n2858), .Z(n710) );
  XNOR U1015 ( .A(n701), .B(n2453), .Z(n847) );
  IV U1016 ( .A(shift_row_out[79]), .Z(n701) );
  NAND U1017 ( .A(n566), .B(shift_row_out[71]), .Z(n844) );
  XOR U1018 ( .A(n849), .B(key[70]), .Z(o[70]) );
  NAND U1019 ( .A(n850), .B(n851), .Z(n849) );
  NAND U1020 ( .A(n556), .B(msg[70]), .Z(n851) );
  AND U1021 ( .A(n852), .B(n853), .Z(n850) );
  NAND U1022 ( .A(n854), .B(n560), .Z(n853) );
  XOR U1023 ( .A(n855), .B(n856), .Z(n854) );
  XNOR U1024 ( .A(n624), .B(n2858), .Z(n856) );
  IV U1025 ( .A(n2452), .Z(n624) );
  XOR U1026 ( .A(n2857), .B(n700), .Z(n855) );
  XOR U1027 ( .A(n787), .B(n2372), .Z(n700) );
  IV U1028 ( .A(n1967), .Z(n787) );
  NANDN U1029 ( .B(n2453), .A(n566), .Z(n852) );
  XOR U1030 ( .A(n857), .B(key[6]), .Z(o[6]) );
  NAND U1031 ( .A(n858), .B(n859), .Z(n857) );
  NAND U1032 ( .A(n556), .B(msg[6]), .Z(n859) );
  AND U1033 ( .A(n860), .B(n861), .Z(n858) );
  NAND U1034 ( .A(n862), .B(n560), .Z(n861) );
  XOR U1035 ( .A(n863), .B(n864), .Z(n862) );
  XNOR U1036 ( .A(n779), .B(n2209), .Z(n864) );
  XOR U1037 ( .A(\b/SBOX[0].sbox/n90 ), .B(n865), .Z(n863) );
  NANDN U1038 ( .B(\b/SBOX[0].sbox/n91 ), .A(n566), .Z(n860) );
  XOR U1039 ( .A(n866), .B(key[69]), .Z(o[69]) );
  NAND U1040 ( .A(n867), .B(n868), .Z(n866) );
  NAND U1041 ( .A(n556), .B(msg[69]), .Z(n868) );
  AND U1042 ( .A(n869), .B(n870), .Z(n867) );
  NAND U1043 ( .A(n871), .B(n560), .Z(n870) );
  XOR U1044 ( .A(n872), .B(n873), .Z(n871) );
  XOR U1045 ( .A(shift_row_out[76]), .B(shift_row_out[68]), .Z(n873) );
  XNOR U1046 ( .A(n720), .B(n711), .Z(n872) );
  XOR U1047 ( .A(n795), .B(n2371), .Z(n711) );
  IV U1048 ( .A(n1966), .Z(n795) );
  IV U1049 ( .A(n2857), .Z(n720) );
  NANDN U1050 ( .B(n2452), .A(n566), .Z(n869) );
  XOR U1051 ( .A(n874), .B(key[68]), .Z(o[68]) );
  NAND U1052 ( .A(n875), .B(n876), .Z(n874) );
  NAND U1053 ( .A(n556), .B(msg[68]), .Z(n876) );
  AND U1054 ( .A(n877), .B(n878), .Z(n875) );
  NAND U1055 ( .A(n879), .B(n560), .Z(n878) );
  XOR U1056 ( .A(n880), .B(n881), .Z(n879) );
  XOR U1057 ( .A(n721), .B(n882), .Z(n881) );
  XNOR U1058 ( .A(shift_row_out[84]), .B(shift_row_out[92]), .Z(n721) );
  XOR U1059 ( .A(shift_row_out[67]), .B(n883), .Z(n880) );
  XOR U1060 ( .A(shift_row_out[76]), .B(shift_row_out[75]), .Z(n883) );
  NAND U1061 ( .A(n566), .B(shift_row_out[68]), .Z(n877) );
  XOR U1062 ( .A(n884), .B(key[67]), .Z(o[67]) );
  NAND U1063 ( .A(n885), .B(n886), .Z(n884) );
  NAND U1064 ( .A(n556), .B(msg[67]), .Z(n886) );
  AND U1065 ( .A(n887), .B(n888), .Z(n885) );
  NAND U1066 ( .A(n889), .B(n560), .Z(n888) );
  XOR U1067 ( .A(n890), .B(n891), .Z(n889) );
  XOR U1068 ( .A(n730), .B(n882), .Z(n891) );
  IV U1069 ( .A(n892), .Z(n882) );
  XNOR U1070 ( .A(shift_row_out[83]), .B(shift_row_out[91]), .Z(n730) );
  XOR U1071 ( .A(shift_row_out[66]), .B(n893), .Z(n890) );
  XOR U1072 ( .A(shift_row_out[75]), .B(shift_row_out[74]), .Z(n893) );
  NAND U1073 ( .A(n566), .B(shift_row_out[67]), .Z(n887) );
  XOR U1074 ( .A(n894), .B(key[66]), .Z(o[66]) );
  NAND U1075 ( .A(n895), .B(n896), .Z(n894) );
  NAND U1076 ( .A(msg[66]), .B(n556), .Z(n896) );
  AND U1077 ( .A(n897), .B(n898), .Z(n895) );
  NAND U1078 ( .A(n899), .B(n560), .Z(n898) );
  XOR U1079 ( .A(n900), .B(n901), .Z(n899) );
  XNOR U1080 ( .A(n2856), .B(n741), .Z(n901) );
  XNOR U1081 ( .A(shift_row_out[82]), .B(shift_row_out[90]), .Z(n741) );
  XOR U1082 ( .A(shift_row_out[74]), .B(n2451), .Z(n900) );
  NAND U1083 ( .A(n566), .B(shift_row_out[66]), .Z(n897) );
  XOR U1084 ( .A(n902), .B(key[65]), .Z(o[65]) );
  NAND U1085 ( .A(n903), .B(n904), .Z(n902) );
  NAND U1086 ( .A(n556), .B(msg[65]), .Z(n904) );
  AND U1087 ( .A(n905), .B(n906), .Z(n903) );
  NAND U1088 ( .A(n907), .B(n560), .Z(n906) );
  XOR U1089 ( .A(n908), .B(n909), .Z(n907) );
  XNOR U1090 ( .A(n751), .B(n892), .Z(n909) );
  XNOR U1091 ( .A(n1965), .B(n2370), .Z(n751) );
  XNOR U1092 ( .A(n2855), .B(n910), .Z(n908) );
  XNOR U1093 ( .A(n683), .B(n2856), .Z(n910) );
  IV U1094 ( .A(n2450), .Z(n683) );
  NANDN U1095 ( .B(n2451), .A(n566), .Z(n905) );
  XOR U1096 ( .A(n911), .B(key[64]), .Z(o[64]) );
  NAND U1097 ( .A(n912), .B(n913), .Z(n911) );
  NAND U1098 ( .A(n556), .B(msg[64]), .Z(n913) );
  AND U1099 ( .A(n914), .B(n915), .Z(n912) );
  NAND U1100 ( .A(n916), .B(n560), .Z(n915) );
  XOR U1101 ( .A(n917), .B(n892), .Z(n916) );
  XOR U1102 ( .A(shift_row_out[71]), .B(shift_row_out[79]), .Z(n892) );
  XOR U1103 ( .A(n2855), .B(n760), .Z(n917) );
  XNOR U1104 ( .A(n1964), .B(n2369), .Z(n760) );
  NANDN U1105 ( .B(n2450), .A(n566), .Z(n914) );
  XOR U1106 ( .A(n918), .B(key[63]), .Z(o[63]) );
  NAND U1107 ( .A(n919), .B(n920), .Z(n918) );
  NAND U1108 ( .A(n556), .B(msg[63]), .Z(n920) );
  AND U1109 ( .A(n921), .B(n922), .Z(n919) );
  NAND U1110 ( .A(n923), .B(n560), .Z(n922) );
  XOR U1111 ( .A(n924), .B(n925), .Z(n923) );
  XOR U1112 ( .A(n2048), .B(n926), .Z(n925) );
  XNOR U1113 ( .A(shift_row_out[39]), .B(n927), .Z(n924) );
  NAND U1114 ( .A(n566), .B(shift_row_out[63]), .Z(n921) );
  XOR U1115 ( .A(n928), .B(key[62]), .Z(o[62]) );
  NAND U1116 ( .A(n929), .B(n930), .Z(n928) );
  NAND U1117 ( .A(n556), .B(msg[62]), .Z(n930) );
  AND U1118 ( .A(n931), .B(n932), .Z(n929) );
  NAND U1119 ( .A(n933), .B(n560), .Z(n932) );
  XOR U1120 ( .A(n934), .B(n935), .Z(n933) );
  XNOR U1121 ( .A(n927), .B(n2128), .Z(n935) );
  XOR U1122 ( .A(n2047), .B(n936), .Z(n934) );
  NANDN U1123 ( .B(n2048), .A(n566), .Z(n931) );
  XOR U1124 ( .A(n937), .B(key[61]), .Z(o[61]) );
  NAND U1125 ( .A(n938), .B(n939), .Z(n937) );
  NAND U1126 ( .A(n556), .B(msg[61]), .Z(n939) );
  AND U1127 ( .A(n940), .B(n941), .Z(n938) );
  NAND U1128 ( .A(n942), .B(n560), .Z(n941) );
  XOR U1129 ( .A(n943), .B(n944), .Z(n942) );
  XOR U1130 ( .A(shift_row_out[60]), .B(shift_row_out[36]), .Z(n944) );
  XOR U1131 ( .A(n2128), .B(n945), .Z(n943) );
  NANDN U1132 ( .B(n2047), .A(n566), .Z(n940) );
  XOR U1133 ( .A(n946), .B(key[60]), .Z(o[60]) );
  NAND U1134 ( .A(n947), .B(n948), .Z(n946) );
  NAND U1135 ( .A(n556), .B(msg[60]), .Z(n948) );
  AND U1136 ( .A(n949), .B(n950), .Z(n947) );
  NAND U1137 ( .A(n951), .B(n560), .Z(n950) );
  XOR U1138 ( .A(n952), .B(n953), .Z(n951) );
  XOR U1139 ( .A(n954), .B(n955), .Z(n953) );
  XOR U1140 ( .A(shift_row_out[35]), .B(n956), .Z(n952) );
  XOR U1141 ( .A(shift_row_out[59]), .B(shift_row_out[36]), .Z(n956) );
  NAND U1142 ( .A(n566), .B(shift_row_out[60]), .Z(n949) );
  XOR U1143 ( .A(n957), .B(key[5]), .Z(o[5]) );
  NAND U1144 ( .A(n958), .B(n959), .Z(n957) );
  NAND U1145 ( .A(n556), .B(msg[5]), .Z(n959) );
  AND U1146 ( .A(n960), .B(n961), .Z(n958) );
  NAND U1147 ( .A(n962), .B(n560), .Z(n961) );
  XOR U1148 ( .A(n963), .B(n964), .Z(n962) );
  XOR U1149 ( .A(shift_row_out[4]), .B(shift_row_out[12]), .Z(n964) );
  XOR U1150 ( .A(n2209), .B(n965), .Z(n963) );
  NANDN U1151 ( .B(\b/SBOX[0].sbox/n90 ), .A(n566), .Z(n960) );
  XOR U1152 ( .A(n966), .B(key[59]), .Z(o[59]) );
  NAND U1153 ( .A(n967), .B(n968), .Z(n966) );
  NAND U1154 ( .A(n556), .B(msg[59]), .Z(n968) );
  AND U1155 ( .A(n969), .B(n970), .Z(n967) );
  NAND U1156 ( .A(n971), .B(n560), .Z(n970) );
  XOR U1157 ( .A(n972), .B(n973), .Z(n971) );
  XOR U1158 ( .A(n954), .B(n974), .Z(n973) );
  XOR U1159 ( .A(shift_row_out[34]), .B(n975), .Z(n972) );
  XOR U1160 ( .A(shift_row_out[58]), .B(shift_row_out[35]), .Z(n975) );
  NAND U1161 ( .A(n566), .B(shift_row_out[59]), .Z(n969) );
  XOR U1162 ( .A(n976), .B(key[58]), .Z(o[58]) );
  NAND U1163 ( .A(n977), .B(n978), .Z(n976) );
  NAND U1164 ( .A(msg[58]), .B(n556), .Z(n978) );
  AND U1165 ( .A(n979), .B(n980), .Z(n977) );
  NAND U1166 ( .A(n981), .B(n560), .Z(n980) );
  XOR U1167 ( .A(n982), .B(n983), .Z(n981) );
  XNOR U1168 ( .A(n2046), .B(n984), .Z(n983) );
  XNOR U1169 ( .A(shift_row_out[34]), .B(n985), .Z(n982) );
  NAND U1170 ( .A(n566), .B(shift_row_out[58]), .Z(n979) );
  XOR U1171 ( .A(n986), .B(key[57]), .Z(o[57]) );
  NAND U1172 ( .A(n987), .B(n988), .Z(n986) );
  NAND U1173 ( .A(n556), .B(msg[57]), .Z(n988) );
  AND U1174 ( .A(n989), .B(n990), .Z(n987) );
  NAND U1175 ( .A(n991), .B(n560), .Z(n990) );
  XOR U1176 ( .A(n992), .B(n993), .Z(n991) );
  XOR U1177 ( .A(n954), .B(n994), .Z(n993) );
  XNOR U1178 ( .A(n2045), .B(n995), .Z(n992) );
  XNOR U1179 ( .A(n985), .B(n2126), .Z(n995) );
  NANDN U1180 ( .B(n2046), .A(n566), .Z(n989) );
  XOR U1181 ( .A(n996), .B(key[56]), .Z(o[56]) );
  NAND U1182 ( .A(n997), .B(n998), .Z(n996) );
  NAND U1183 ( .A(n556), .B(msg[56]), .Z(n998) );
  AND U1184 ( .A(n999), .B(n1000), .Z(n997) );
  NAND U1185 ( .A(n1001), .B(n560), .Z(n1000) );
  XNOR U1186 ( .A(n1002), .B(n1003), .Z(n1001) );
  XOR U1187 ( .A(n2126), .B(n954), .Z(n1002) );
  XNOR U1188 ( .A(shift_row_out[39]), .B(shift_row_out[63]), .Z(n954) );
  NANDN U1189 ( .B(n2045), .A(n566), .Z(n999) );
  XOR U1190 ( .A(n1004), .B(key[55]), .Z(o[55]) );
  NAND U1191 ( .A(n1005), .B(n1006), .Z(n1004) );
  NAND U1192 ( .A(n556), .B(msg[55]), .Z(n1006) );
  AND U1193 ( .A(n1007), .B(n1008), .Z(n1005) );
  NAND U1194 ( .A(n1009), .B(n560), .Z(n1008) );
  XOR U1195 ( .A(n1010), .B(n1011), .Z(n1009) );
  XNOR U1196 ( .A(shift_row_out[39]), .B(n1012), .Z(n1011) );
  XOR U1197 ( .A(shift_row_out[63]), .B(shift_row_out[47]), .Z(n1010) );
  NAND U1198 ( .A(n566), .B(shift_row_out[55]), .Z(n1007) );
  XOR U1199 ( .A(n1013), .B(key[54]), .Z(o[54]) );
  NAND U1200 ( .A(n1014), .B(n1015), .Z(n1013) );
  NAND U1201 ( .A(n556), .B(msg[54]), .Z(n1015) );
  AND U1202 ( .A(n1016), .B(n1017), .Z(n1014) );
  NAND U1203 ( .A(n1018), .B(n560), .Z(n1017) );
  XOR U1204 ( .A(n1019), .B(n1020), .Z(n1018) );
  XNOR U1205 ( .A(n2534), .B(n927), .Z(n1020) );
  XNOR U1206 ( .A(n2048), .B(n1021), .Z(n1019) );
  NANDN U1207 ( .B(n2939), .A(n566), .Z(n1016) );
  XOR U1208 ( .A(n1022), .B(key[53]), .Z(o[53]) );
  NAND U1209 ( .A(n1023), .B(n1024), .Z(n1022) );
  NAND U1210 ( .A(n556), .B(msg[53]), .Z(n1024) );
  AND U1211 ( .A(n1025), .B(n1026), .Z(n1023) );
  NAND U1212 ( .A(n1027), .B(n560), .Z(n1026) );
  XOR U1213 ( .A(n1028), .B(n1029), .Z(n1027) );
  XNOR U1214 ( .A(n1030), .B(n2128), .Z(n1029) );
  XOR U1215 ( .A(n2047), .B(n1031), .Z(n1028) );
  NANDN U1216 ( .B(n2938), .A(n566), .Z(n1025) );
  XOR U1217 ( .A(n1032), .B(key[52]), .Z(o[52]) );
  NAND U1218 ( .A(n1033), .B(n1034), .Z(n1032) );
  NAND U1219 ( .A(n556), .B(msg[52]), .Z(n1034) );
  AND U1220 ( .A(n1035), .B(n1036), .Z(n1033) );
  NAND U1221 ( .A(n1037), .B(n560), .Z(n1036) );
  XOR U1222 ( .A(n1038), .B(n1039), .Z(n1037) );
  XNOR U1223 ( .A(n1040), .B(n1041), .Z(n1039) );
  XOR U1224 ( .A(shift_row_out[36]), .B(n1042), .Z(n1038) );
  XOR U1225 ( .A(shift_row_out[60]), .B(shift_row_out[44]), .Z(n1042) );
  NAND U1226 ( .A(n566), .B(shift_row_out[52]), .Z(n1035) );
  XOR U1227 ( .A(n1043), .B(key[51]), .Z(o[51]) );
  NAND U1228 ( .A(n1044), .B(n1045), .Z(n1043) );
  NAND U1229 ( .A(n556), .B(msg[51]), .Z(n1045) );
  AND U1230 ( .A(n1046), .B(n1047), .Z(n1044) );
  NAND U1231 ( .A(n1048), .B(n560), .Z(n1047) );
  XOR U1232 ( .A(n1049), .B(n1050), .Z(n1048) );
  XNOR U1233 ( .A(n1041), .B(n1051), .Z(n1050) );
  XOR U1234 ( .A(shift_row_out[35]), .B(n1052), .Z(n1049) );
  XOR U1235 ( .A(shift_row_out[59]), .B(shift_row_out[43]), .Z(n1052) );
  NAND U1236 ( .A(n566), .B(shift_row_out[51]), .Z(n1046) );
  XOR U1237 ( .A(n1053), .B(key[50]), .Z(o[50]) );
  NAND U1238 ( .A(n1054), .B(n1055), .Z(n1053) );
  NAND U1239 ( .A(msg[50]), .B(n556), .Z(n1055) );
  AND U1240 ( .A(n1056), .B(n1057), .Z(n1054) );
  NAND U1241 ( .A(n1058), .B(n560), .Z(n1057) );
  XOR U1242 ( .A(n1059), .B(n1060), .Z(n1058) );
  XOR U1243 ( .A(shift_row_out[34]), .B(n1061), .Z(n1060) );
  XOR U1244 ( .A(shift_row_out[58]), .B(shift_row_out[42]), .Z(n1059) );
  NAND U1245 ( .A(n566), .B(shift_row_out[50]), .Z(n1056) );
  XOR U1246 ( .A(n1062), .B(key[4]), .Z(o[4]) );
  NAND U1247 ( .A(n1063), .B(n1064), .Z(n1062) );
  NAND U1248 ( .A(n556), .B(msg[4]), .Z(n1064) );
  AND U1249 ( .A(n1065), .B(n1066), .Z(n1063) );
  NAND U1250 ( .A(n1067), .B(n560), .Z(n1066) );
  XOR U1251 ( .A(n1068), .B(n1069), .Z(n1067) );
  XOR U1252 ( .A(n1070), .B(n1071), .Z(n1069) );
  XOR U1253 ( .A(shift_row_out[11]), .B(n1072), .Z(n1068) );
  XOR U1254 ( .A(shift_row_out[3]), .B(shift_row_out[12]), .Z(n1072) );
  NAND U1255 ( .A(n566), .B(shift_row_out[4]), .Z(n1065) );
  XOR U1256 ( .A(n1073), .B(key[49]), .Z(o[49]) );
  NAND U1257 ( .A(n1074), .B(n1075), .Z(n1073) );
  NAND U1258 ( .A(n556), .B(msg[49]), .Z(n1075) );
  AND U1259 ( .A(n1076), .B(n1077), .Z(n1074) );
  NAND U1260 ( .A(n1078), .B(n560), .Z(n1077) );
  XOR U1261 ( .A(n1079), .B(n1080), .Z(n1078) );
  XNOR U1262 ( .A(n1081), .B(n1082), .Z(n1080) );
  XNOR U1263 ( .A(n2046), .B(n1083), .Z(n1079) );
  XNOR U1264 ( .A(n2532), .B(n985), .Z(n1083) );
  NANDN U1265 ( .B(n2937), .A(n566), .Z(n1076) );
  XOR U1266 ( .A(n1084), .B(key[48]), .Z(o[48]) );
  NAND U1267 ( .A(n1085), .B(n1086), .Z(n1084) );
  NAND U1268 ( .A(n556), .B(msg[48]), .Z(n1086) );
  AND U1269 ( .A(n1087), .B(n1088), .Z(n1085) );
  NAND U1270 ( .A(n1089), .B(n560), .Z(n1088) );
  XOR U1271 ( .A(n1090), .B(n1091), .Z(n1089) );
  XNOR U1272 ( .A(n1092), .B(n2126), .Z(n1091) );
  XNOR U1273 ( .A(n2045), .B(n1041), .Z(n1090) );
  NANDN U1274 ( .B(n2936), .A(n566), .Z(n1087) );
  XOR U1275 ( .A(n1093), .B(key[47]), .Z(o[47]) );
  NAND U1276 ( .A(n1094), .B(n1095), .Z(n1093) );
  NAND U1277 ( .A(n556), .B(msg[47]), .Z(n1095) );
  AND U1278 ( .A(n1096), .B(n1097), .Z(n1094) );
  NAND U1279 ( .A(n1098), .B(n560), .Z(n1097) );
  XOR U1280 ( .A(n1041), .B(n1099), .Z(n1098) );
  XNOR U1281 ( .A(shift_row_out[39]), .B(n936), .Z(n1099) );
  XNOR U1282 ( .A(n2939), .B(n2534), .Z(n936) );
  IV U1283 ( .A(n1081), .Z(n1041) );
  NAND U1284 ( .A(shift_row_out[47]), .B(n566), .Z(n1096) );
  XOR U1285 ( .A(n1100), .B(key[46]), .Z(o[46]) );
  NAND U1286 ( .A(n1101), .B(n1102), .Z(n1100) );
  NAND U1287 ( .A(n556), .B(msg[46]), .Z(n1102) );
  AND U1288 ( .A(n1103), .B(n1104), .Z(n1101) );
  NAND U1289 ( .A(n1105), .B(n560), .Z(n1104) );
  XOR U1290 ( .A(n2129), .B(n945), .Z(n1106) );
  XNOR U1291 ( .A(n2938), .B(n2533), .Z(n945) );
  NANDN U1292 ( .B(n2534), .A(n566), .Z(n1103) );
  XOR U1293 ( .A(n1107), .B(key[45]), .Z(o[45]) );
  NAND U1294 ( .A(n1108), .B(n1109), .Z(n1107) );
  NAND U1295 ( .A(n556), .B(msg[45]), .Z(n1109) );
  AND U1296 ( .A(n1110), .B(n1111), .Z(n1108) );
  NAND U1297 ( .A(n1112), .B(n560), .Z(n1111) );
  XOR U1298 ( .A(n1113), .B(n1021), .Z(n1112) );
  XOR U1299 ( .A(n2128), .B(n955), .Z(n1113) );
  XNOR U1300 ( .A(shift_row_out[44]), .B(shift_row_out[52]), .Z(n955) );
  NANDN U1301 ( .B(n2533), .A(n566), .Z(n1110) );
  XOR U1302 ( .A(n1114), .B(key[44]), .Z(o[44]) );
  NAND U1303 ( .A(n1115), .B(n1116), .Z(n1114) );
  NAND U1304 ( .A(n556), .B(msg[44]), .Z(n1116) );
  AND U1305 ( .A(n1117), .B(n1118), .Z(n1115) );
  NAND U1306 ( .A(n1119), .B(n560), .Z(n1118) );
  XOR U1307 ( .A(n1120), .B(n1121), .Z(n1119) );
  XOR U1308 ( .A(n974), .B(n1031), .Z(n1121) );
  XNOR U1309 ( .A(shift_row_out[43]), .B(shift_row_out[51]), .Z(n974) );
  XOR U1310 ( .A(shift_row_out[36]), .B(n926), .Z(n1120) );
  NAND U1311 ( .A(n566), .B(shift_row_out[44]), .Z(n1117) );
  XOR U1312 ( .A(n1122), .B(key[43]), .Z(o[43]) );
  NAND U1313 ( .A(n1123), .B(n1124), .Z(n1122) );
  NAND U1314 ( .A(n556), .B(msg[43]), .Z(n1124) );
  AND U1315 ( .A(n1125), .B(n1126), .Z(n1123) );
  NAND U1316 ( .A(n1127), .B(n560), .Z(n1126) );
  XOR U1317 ( .A(n1128), .B(n1129), .Z(n1127) );
  XOR U1318 ( .A(n984), .B(n1040), .Z(n1129) );
  XNOR U1319 ( .A(shift_row_out[42]), .B(shift_row_out[50]), .Z(n984) );
  XOR U1320 ( .A(shift_row_out[35]), .B(n926), .Z(n1128) );
  NAND U1321 ( .A(n566), .B(shift_row_out[43]), .Z(n1125) );
  XOR U1322 ( .A(n1130), .B(key[42]), .Z(o[42]) );
  NAND U1323 ( .A(n1131), .B(n1132), .Z(n1130) );
  NAND U1324 ( .A(msg[42]), .B(n556), .Z(n1132) );
  AND U1325 ( .A(n1133), .B(n1134), .Z(n1131) );
  NAND U1326 ( .A(n1135), .B(n560), .Z(n1134) );
  XNOR U1327 ( .A(n1051), .B(n1136), .Z(n1135) );
  XNOR U1328 ( .A(shift_row_out[34]), .B(n994), .Z(n1136) );
  XNOR U1329 ( .A(n2937), .B(n2532), .Z(n994) );
  NAND U1330 ( .A(n566), .B(shift_row_out[42]), .Z(n1133) );
  XOR U1331 ( .A(n1137), .B(key[41]), .Z(o[41]) );
  NAND U1332 ( .A(n1138), .B(n1139), .Z(n1137) );
  NAND U1333 ( .A(n556), .B(msg[41]), .Z(n1139) );
  AND U1334 ( .A(n1140), .B(n1141), .Z(n1138) );
  NAND U1335 ( .A(n1142), .B(n560), .Z(n1141) );
  XOR U1336 ( .A(n1143), .B(n1144), .Z(n1142) );
  XNOR U1337 ( .A(n1003), .B(n1061), .Z(n1144) );
  XNOR U1338 ( .A(n2936), .B(n2531), .Z(n1003) );
  XNOR U1339 ( .A(n2127), .B(n926), .Z(n1143) );
  NANDN U1340 ( .B(n2532), .A(n566), .Z(n1140) );
  XOR U1341 ( .A(n1145), .B(key[40]), .Z(o[40]) );
  NAND U1342 ( .A(n1146), .B(n1147), .Z(n1145) );
  NAND U1343 ( .A(n556), .B(msg[40]), .Z(n1147) );
  AND U1344 ( .A(n1148), .B(n1149), .Z(n1146) );
  NAND U1345 ( .A(n1150), .B(n560), .Z(n1149) );
  XOR U1346 ( .A(n1151), .B(n1082), .Z(n1150) );
  XNOR U1347 ( .A(n2126), .B(n926), .Z(n1151) );
  XOR U1348 ( .A(shift_row_out[47]), .B(shift_row_out[55]), .Z(n926) );
  NANDN U1349 ( .B(n2531), .A(n566), .Z(n1148) );
  XOR U1350 ( .A(n1152), .B(key[3]), .Z(o[3]) );
  NAND U1351 ( .A(n1153), .B(n1154), .Z(n1152) );
  NAND U1352 ( .A(n556), .B(msg[3]), .Z(n1154) );
  AND U1353 ( .A(n1155), .B(n1156), .Z(n1153) );
  NAND U1354 ( .A(n1157), .B(n560), .Z(n1156) );
  XOR U1355 ( .A(n1158), .B(n1159), .Z(n1157) );
  XOR U1356 ( .A(n1070), .B(n1160), .Z(n1159) );
  XOR U1357 ( .A(shift_row_out[10]), .B(n1161), .Z(n1158) );
  XOR U1358 ( .A(shift_row_out[2]), .B(shift_row_out[11]), .Z(n1161) );
  NAND U1359 ( .A(n566), .B(shift_row_out[3]), .Z(n1155) );
  XOR U1360 ( .A(n1162), .B(key[39]), .Z(o[39]) );
  NAND U1361 ( .A(n1163), .B(n1164), .Z(n1162) );
  NAND U1362 ( .A(n556), .B(msg[39]), .Z(n1164) );
  AND U1363 ( .A(n1165), .B(n1166), .Z(n1163) );
  NAND U1364 ( .A(n1167), .B(n560), .Z(n1166) );
  XOR U1365 ( .A(n1168), .B(n1169), .Z(n1167) );
  XOR U1366 ( .A(n927), .B(n1081), .Z(n1169) );
  XNOR U1367 ( .A(shift_row_out[55]), .B(shift_row_out[63]), .Z(n1081) );
  IV U1368 ( .A(n2129), .Z(n927) );
  XOR U1369 ( .A(shift_row_out[47]), .B(n2534), .Z(n1168) );
  NAND U1370 ( .A(n566), .B(shift_row_out[39]), .Z(n1165) );
  XOR U1371 ( .A(n1170), .B(key[38]), .Z(o[38]) );
  NAND U1372 ( .A(n1171), .B(n1172), .Z(n1170) );
  NAND U1373 ( .A(n556), .B(msg[38]), .Z(n1172) );
  AND U1374 ( .A(n1173), .B(n1174), .Z(n1171) );
  NAND U1375 ( .A(n1175), .B(n560), .Z(n1174) );
  XOR U1376 ( .A(n1176), .B(n1177), .Z(n1175) );
  XNOR U1377 ( .A(n2534), .B(n1030), .Z(n1177) );
  XOR U1378 ( .A(n2128), .B(n1012), .Z(n1176) );
  NANDN U1379 ( .B(n2129), .A(n566), .Z(n1173) );
  XOR U1380 ( .A(n1178), .B(key[37]), .Z(o[37]) );
  NAND U1381 ( .A(n1179), .B(n1180), .Z(n1178) );
  NAND U1382 ( .A(n556), .B(msg[37]), .Z(n1180) );
  AND U1383 ( .A(n1181), .B(n1182), .Z(n1179) );
  NAND U1384 ( .A(n1183), .B(n560), .Z(n1182) );
  XOR U1385 ( .A(n1184), .B(n1185), .Z(n1183) );
  XOR U1386 ( .A(shift_row_out[44]), .B(shift_row_out[36]), .Z(n1185) );
  XOR U1387 ( .A(n1030), .B(n1021), .Z(n1184) );
  IV U1388 ( .A(n2533), .Z(n1030) );
  NANDN U1389 ( .B(n2128), .A(n566), .Z(n1181) );
  XOR U1390 ( .A(n1186), .B(key[36]), .Z(o[36]) );
  NAND U1391 ( .A(n1187), .B(n1188), .Z(n1186) );
  NAND U1392 ( .A(n556), .B(msg[36]), .Z(n1188) );
  AND U1393 ( .A(n1189), .B(n1190), .Z(n1187) );
  NAND U1394 ( .A(n1191), .B(n560), .Z(n1190) );
  XOR U1395 ( .A(n1192), .B(n1193), .Z(n1191) );
  XOR U1396 ( .A(n1031), .B(n1194), .Z(n1193) );
  XNOR U1397 ( .A(shift_row_out[52]), .B(shift_row_out[60]), .Z(n1031) );
  XOR U1398 ( .A(shift_row_out[35]), .B(n1195), .Z(n1192) );
  XOR U1399 ( .A(shift_row_out[44]), .B(shift_row_out[43]), .Z(n1195) );
  NAND U1400 ( .A(n566), .B(shift_row_out[36]), .Z(n1189) );
  XOR U1401 ( .A(n1196), .B(key[35]), .Z(o[35]) );
  NAND U1402 ( .A(n1197), .B(n1198), .Z(n1196) );
  NAND U1403 ( .A(n556), .B(msg[35]), .Z(n1198) );
  AND U1404 ( .A(n1199), .B(n1200), .Z(n1197) );
  NAND U1405 ( .A(n1201), .B(n560), .Z(n1200) );
  XOR U1406 ( .A(n1202), .B(n1203), .Z(n1201) );
  XOR U1407 ( .A(n1040), .B(n1194), .Z(n1203) );
  XNOR U1408 ( .A(shift_row_out[51]), .B(shift_row_out[59]), .Z(n1040) );
  XOR U1409 ( .A(shift_row_out[34]), .B(n1204), .Z(n1202) );
  XOR U1410 ( .A(shift_row_out[43]), .B(shift_row_out[42]), .Z(n1204) );
  NAND U1411 ( .A(n566), .B(shift_row_out[35]), .Z(n1199) );
  XOR U1412 ( .A(n1205), .B(key[34]), .Z(o[34]) );
  NAND U1413 ( .A(n1206), .B(n1207), .Z(n1205) );
  NAND U1414 ( .A(msg[34]), .B(n556), .Z(n1207) );
  AND U1415 ( .A(n1208), .B(n1209), .Z(n1206) );
  NAND U1416 ( .A(n1210), .B(n560), .Z(n1209) );
  XOR U1417 ( .A(n1211), .B(n1212), .Z(n1210) );
  XOR U1418 ( .A(n985), .B(n1051), .Z(n1212) );
  XNOR U1419 ( .A(shift_row_out[50]), .B(shift_row_out[58]), .Z(n1051) );
  IV U1420 ( .A(n2127), .Z(n985) );
  XOR U1421 ( .A(shift_row_out[42]), .B(n2532), .Z(n1211) );
  NAND U1422 ( .A(n566), .B(shift_row_out[34]), .Z(n1208) );
  XOR U1423 ( .A(n1213), .B(key[33]), .Z(o[33]) );
  NAND U1424 ( .A(n1214), .B(n1215), .Z(n1213) );
  NAND U1425 ( .A(n556), .B(msg[33]), .Z(n1215) );
  AND U1426 ( .A(n1216), .B(n1217), .Z(n1214) );
  NAND U1427 ( .A(n1218), .B(n560), .Z(n1217) );
  XOR U1428 ( .A(n1219), .B(n1220), .Z(n1218) );
  XNOR U1429 ( .A(n1061), .B(n1194), .Z(n1220) );
  IV U1430 ( .A(n1221), .Z(n1194) );
  XNOR U1431 ( .A(n2126), .B(n1222), .Z(n1219) );
  XNOR U1432 ( .A(n2532), .B(n1092), .Z(n1222) );
  NANDN U1433 ( .B(n2127), .A(n566), .Z(n1216) );
  XOR U1434 ( .A(n1223), .B(key[32]), .Z(o[32]) );
  NAND U1435 ( .A(n1224), .B(n1225), .Z(n1223) );
  NAND U1436 ( .A(n556), .B(msg[32]), .Z(n1225) );
  AND U1437 ( .A(n1226), .B(n1227), .Z(n1224) );
  NAND U1438 ( .A(n1228), .B(n560), .Z(n1227) );
  XOR U1439 ( .A(n1229), .B(n1221), .Z(n1228) );
  XOR U1440 ( .A(shift_row_out[39]), .B(shift_row_out[47]), .Z(n1221) );
  XOR U1441 ( .A(n1092), .B(n1082), .Z(n1229) );
  IV U1442 ( .A(n2531), .Z(n1092) );
  NANDN U1443 ( .B(n2126), .A(n566), .Z(n1226) );
  XOR U1444 ( .A(n1230), .B(key[31]), .Z(o[31]) );
  NAND U1445 ( .A(n1231), .B(n1232), .Z(n1230) );
  NAND U1446 ( .A(n556), .B(msg[31]), .Z(n1232) );
  AND U1447 ( .A(n1233), .B(n1234), .Z(n1231) );
  NAND U1448 ( .A(n1235), .B(n560), .Z(n1234) );
  XOR U1449 ( .A(n1236), .B(n1237), .Z(n1235) );
  XNOR U1450 ( .A(shift_row_out[15]), .B(n1238), .Z(n1237) );
  XOR U1451 ( .A(shift_row_out[7]), .B(shift_row_out[23]), .Z(n1236) );
  NAND U1452 ( .A(n566), .B(shift_row_out[31]), .Z(n1233) );
  XOR U1453 ( .A(n1239), .B(key[30]), .Z(o[30]) );
  NAND U1454 ( .A(n1240), .B(n1241), .Z(n1239) );
  NAND U1455 ( .A(n556), .B(msg[30]), .Z(n1241) );
  AND U1456 ( .A(n1242), .B(n1243), .Z(n1240) );
  NAND U1457 ( .A(n1244), .B(n560), .Z(n1243) );
  XOR U1458 ( .A(n1245), .B(n1246), .Z(n1244) );
  XNOR U1459 ( .A(n779), .B(n2615), .Z(n1246) );
  XOR U1460 ( .A(\b/SBOX[0].sbox/n91 ), .B(n1247), .Z(n1245) );
  NANDN U1461 ( .B(n3020), .A(n566), .Z(n1242) );
  XOR U1462 ( .A(n1248), .B(key[2]), .Z(o[2]) );
  NAND U1463 ( .A(n1249), .B(n1250), .Z(n1248) );
  NAND U1464 ( .A(msg[2]), .B(n556), .Z(n1250) );
  AND U1465 ( .A(n1251), .B(n1252), .Z(n1249) );
  NAND U1466 ( .A(n1253), .B(n560), .Z(n1252) );
  XNOR U1467 ( .A(n1254), .B(n1255), .Z(n1253) );
  XNOR U1468 ( .A(shift_row_out[10]), .B(n1256), .Z(n1255) );
  NAND U1469 ( .A(n566), .B(shift_row_out[2]), .Z(n1251) );
  XOR U1470 ( .A(n1257), .B(key[29]), .Z(o[29]) );
  NAND U1471 ( .A(n1258), .B(n1259), .Z(n1257) );
  NAND U1472 ( .A(n556), .B(msg[29]), .Z(n1259) );
  AND U1473 ( .A(n1260), .B(n1261), .Z(n1258) );
  NAND U1474 ( .A(n1262), .B(n560), .Z(n1261) );
  XOR U1475 ( .A(n1263), .B(n1264), .Z(n1262) );
  XNOR U1476 ( .A(n1265), .B(n2614), .Z(n1264) );
  XOR U1477 ( .A(\b/SBOX[0].sbox/n90 ), .B(n1266), .Z(n1263) );
  NANDN U1478 ( .B(n3019), .A(n566), .Z(n1260) );
  XOR U1479 ( .A(n1267), .B(key[28]), .Z(o[28]) );
  NAND U1480 ( .A(n1268), .B(n1269), .Z(n1267) );
  NAND U1481 ( .A(n556), .B(msg[28]), .Z(n1269) );
  AND U1482 ( .A(n1270), .B(n1271), .Z(n1268) );
  NAND U1483 ( .A(n1272), .B(n560), .Z(n1271) );
  XOR U1484 ( .A(n1273), .B(n1274), .Z(n1272) );
  XNOR U1485 ( .A(n1275), .B(n1276), .Z(n1274) );
  XOR U1486 ( .A(shift_row_out[12]), .B(n1277), .Z(n1273) );
  XOR U1487 ( .A(shift_row_out[4]), .B(shift_row_out[20]), .Z(n1277) );
  NAND U1488 ( .A(n566), .B(shift_row_out[28]), .Z(n1270) );
  XOR U1489 ( .A(n1278), .B(key[27]), .Z(o[27]) );
  NAND U1490 ( .A(n1279), .B(n1280), .Z(n1278) );
  NAND U1491 ( .A(n556), .B(msg[27]), .Z(n1280) );
  AND U1492 ( .A(n1281), .B(n1282), .Z(n1279) );
  NAND U1493 ( .A(n1283), .B(n560), .Z(n1282) );
  XOR U1494 ( .A(n1284), .B(n1285), .Z(n1283) );
  XNOR U1495 ( .A(n1276), .B(n1286), .Z(n1285) );
  XOR U1496 ( .A(shift_row_out[11]), .B(n1287), .Z(n1284) );
  XOR U1497 ( .A(shift_row_out[3]), .B(shift_row_out[19]), .Z(n1287) );
  NAND U1498 ( .A(n566), .B(shift_row_out[27]), .Z(n1281) );
  XOR U1499 ( .A(n1288), .B(key[26]), .Z(o[26]) );
  NAND U1500 ( .A(n1289), .B(n1290), .Z(n1288) );
  NAND U1501 ( .A(msg[26]), .B(n556), .Z(n1290) );
  AND U1502 ( .A(n1291), .B(n1292), .Z(n1289) );
  NAND U1503 ( .A(n1293), .B(n560), .Z(n1292) );
  XOR U1504 ( .A(n1294), .B(n1295), .Z(n1293) );
  XNOR U1505 ( .A(shift_row_out[10]), .B(n563), .Z(n1295) );
  XNOR U1506 ( .A(\b/SBOX[0].sbox/n89 ), .B(n3018), .Z(n563) );
  XOR U1507 ( .A(shift_row_out[2]), .B(shift_row_out[18]), .Z(n1294) );
  NAND U1508 ( .A(n566), .B(shift_row_out[26]), .Z(n1291) );
  XOR U1509 ( .A(n1296), .B(key[25]), .Z(o[25]) );
  NAND U1510 ( .A(n1297), .B(n1298), .Z(n1296) );
  NAND U1511 ( .A(n556), .B(msg[25]), .Z(n1298) );
  AND U1512 ( .A(n1299), .B(n1300), .Z(n1297) );
  NAND U1513 ( .A(n1301), .B(n560), .Z(n1300) );
  XOR U1514 ( .A(n1302), .B(n1303), .Z(n1301) );
  XOR U1515 ( .A(n1254), .B(n1304), .Z(n1303) );
  XNOR U1516 ( .A(\b/SBOX[0].sbox/n89 ), .B(n2208), .Z(n1254) );
  XNOR U1517 ( .A(\b/SBOX[0].sbox/n88 ), .B(n1305), .Z(n1302) );
  XOR U1518 ( .A(n3017), .B(n2613), .Z(n1305) );
  NANDN U1519 ( .B(n3018), .A(n566), .Z(n1299) );
  XOR U1520 ( .A(n1306), .B(key[24]), .Z(o[24]) );
  NAND U1521 ( .A(n1307), .B(n1308), .Z(n1306) );
  NAND U1522 ( .A(n556), .B(msg[24]), .Z(n1308) );
  AND U1523 ( .A(n1309), .B(n1310), .Z(n1307) );
  NAND U1524 ( .A(n1311), .B(n560), .Z(n1310) );
  XNOR U1525 ( .A(n1312), .B(n1304), .Z(n1311) );
  XOR U1526 ( .A(\b/SBOX[0].sbox/n88 ), .B(n565), .Z(n1312) );
  XNOR U1527 ( .A(n2612), .B(n2207), .Z(n565) );
  NANDN U1528 ( .B(n3017), .A(n566), .Z(n1309) );
  XOR U1529 ( .A(n1313), .B(key[23]), .Z(o[23]) );
  NAND U1530 ( .A(n1314), .B(n1315), .Z(n1313) );
  NAND U1531 ( .A(n556), .B(msg[23]), .Z(n1315) );
  AND U1532 ( .A(n1316), .B(n1317), .Z(n1314) );
  NAND U1533 ( .A(n1318), .B(n560), .Z(n1317) );
  XOR U1534 ( .A(n1276), .B(n1319), .Z(n1318) );
  XNOR U1535 ( .A(shift_row_out[15]), .B(n865), .Z(n1319) );
  XNOR U1536 ( .A(n2615), .B(n3020), .Z(n865) );
  NAND U1537 ( .A(shift_row_out[23]), .B(n566), .Z(n1316) );
  XOR U1538 ( .A(n1320), .B(key[22]), .Z(o[22]) );
  NAND U1539 ( .A(n1321), .B(n1322), .Z(n1320) );
  NAND U1540 ( .A(n556), .B(msg[22]), .Z(n1322) );
  AND U1541 ( .A(n1323), .B(n1324), .Z(n1321) );
  NAND U1542 ( .A(n1325), .B(n560), .Z(n1324) );
  XNOR U1543 ( .A(n1326), .B(n1238), .Z(n1325) );
  XOR U1544 ( .A(n2210), .B(n965), .Z(n1326) );
  XNOR U1545 ( .A(n2614), .B(n3019), .Z(n965) );
  NANDN U1546 ( .B(n2615), .A(n566), .Z(n1323) );
  XOR U1547 ( .A(n1327), .B(key[21]), .Z(o[21]) );
  NAND U1548 ( .A(n1328), .B(n1329), .Z(n1327) );
  NAND U1549 ( .A(n556), .B(msg[21]), .Z(n1329) );
  AND U1550 ( .A(n1330), .B(n1331), .Z(n1328) );
  NAND U1551 ( .A(n1332), .B(n560), .Z(n1331) );
  XNOR U1552 ( .A(n1333), .B(n1247), .Z(n1332) );
  XOR U1553 ( .A(n2209), .B(n1071), .Z(n1333) );
  XNOR U1554 ( .A(shift_row_out[20]), .B(shift_row_out[28]), .Z(n1071) );
  NANDN U1555 ( .B(n2614), .A(n566), .Z(n1330) );
  XOR U1556 ( .A(n1334), .B(key[20]), .Z(o[20]) );
  NAND U1557 ( .A(n1335), .B(n1336), .Z(n1334) );
  NAND U1558 ( .A(n556), .B(msg[20]), .Z(n1336) );
  AND U1559 ( .A(n1337), .B(n1338), .Z(n1335) );
  NAND U1560 ( .A(n1339), .B(n560), .Z(n1338) );
  XOR U1561 ( .A(n1340), .B(n1341), .Z(n1339) );
  XOR U1562 ( .A(n1160), .B(n1266), .Z(n1341) );
  XNOR U1563 ( .A(shift_row_out[19]), .B(shift_row_out[27]), .Z(n1160) );
  XNOR U1564 ( .A(shift_row_out[12]), .B(n1342), .Z(n1340) );
  NAND U1565 ( .A(n566), .B(shift_row_out[20]), .Z(n1337) );
  XOR U1566 ( .A(n1343), .B(key[1]), .Z(o[1]) );
  NAND U1567 ( .A(n1344), .B(n1345), .Z(n1343) );
  NAND U1568 ( .A(n556), .B(msg[1]), .Z(n1345) );
  AND U1569 ( .A(n1346), .B(n1347), .Z(n1344) );
  NAND U1570 ( .A(n1348), .B(n560), .Z(n1347) );
  XOR U1571 ( .A(n1349), .B(n1350), .Z(n1348) );
  XOR U1572 ( .A(n1070), .B(n1351), .Z(n1350) );
  XNOR U1573 ( .A(\b/SBOX[0].sbox/n88 ), .B(n1352), .Z(n1349) );
  XNOR U1574 ( .A(n2207), .B(n1353), .Z(n1352) );
  NANDN U1575 ( .B(\b/SBOX[0].sbox/n89 ), .A(n566), .Z(n1346) );
  XOR U1576 ( .A(n1354), .B(key[19]), .Z(o[19]) );
  NAND U1577 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1578 ( .A(n556), .B(msg[19]), .Z(n1356) );
  AND U1579 ( .A(n1357), .B(n1358), .Z(n1355) );
  NAND U1580 ( .A(n1359), .B(n560), .Z(n1358) );
  XOR U1581 ( .A(n1360), .B(n1361), .Z(n1359) );
  XOR U1582 ( .A(n1256), .B(n1275), .Z(n1361) );
  XNOR U1583 ( .A(shift_row_out[18]), .B(shift_row_out[26]), .Z(n1256) );
  XNOR U1584 ( .A(shift_row_out[11]), .B(n1342), .Z(n1360) );
  NAND U1585 ( .A(n566), .B(shift_row_out[19]), .Z(n1357) );
  XOR U1586 ( .A(n1362), .B(key[18]), .Z(o[18]) );
  NAND U1587 ( .A(n1363), .B(n1364), .Z(n1362) );
  NAND U1588 ( .A(msg[18]), .B(n556), .Z(n1364) );
  AND U1589 ( .A(n1365), .B(n1366), .Z(n1363) );
  NAND U1590 ( .A(n1367), .B(n560), .Z(n1366) );
  XOR U1591 ( .A(n1368), .B(n1369), .Z(n1367) );
  XOR U1592 ( .A(shift_row_out[10]), .B(n3018), .Z(n1368) );
  NAND U1593 ( .A(n566), .B(shift_row_out[18]), .Z(n1365) );
  XOR U1594 ( .A(n1370), .B(key[17]), .Z(o[17]) );
  NAND U1595 ( .A(n1371), .B(n1372), .Z(n1370) );
  NAND U1596 ( .A(n556), .B(msg[17]), .Z(n1372) );
  AND U1597 ( .A(n1373), .B(n1374), .Z(n1371) );
  NAND U1598 ( .A(n1375), .B(n560), .Z(n1374) );
  XOR U1599 ( .A(n1376), .B(n1377), .Z(n1375) );
  XNOR U1600 ( .A(n778), .B(n1351), .Z(n1377) );
  XNOR U1601 ( .A(n3018), .B(n2208), .Z(n1351) );
  XOR U1602 ( .A(\b/SBOX[0].sbox/n89 ), .B(n672), .Z(n1376) );
  XNOR U1603 ( .A(n2612), .B(n3017), .Z(n672) );
  NANDN U1604 ( .B(n2613), .A(n566), .Z(n1373) );
  XOR U1605 ( .A(n1378), .B(key[16]), .Z(o[16]) );
  NAND U1606 ( .A(n1379), .B(n1380), .Z(n1378) );
  NAND U1607 ( .A(n556), .B(msg[16]), .Z(n1380) );
  AND U1608 ( .A(n1381), .B(n1382), .Z(n1379) );
  NAND U1609 ( .A(n1383), .B(n560), .Z(n1382) );
  XNOR U1610 ( .A(n1384), .B(n1385), .Z(n1383) );
  XOR U1611 ( .A(\b/SBOX[0].sbox/n88 ), .B(n1342), .Z(n1384) );
  IV U1612 ( .A(n778), .Z(n1342) );
  XOR U1613 ( .A(shift_row_out[23]), .B(shift_row_out[31]), .Z(n778) );
  NANDN U1614 ( .B(n2612), .A(n566), .Z(n1381) );
  XOR U1615 ( .A(n1386), .B(key[15]), .Z(o[15]) );
  NAND U1616 ( .A(n1387), .B(n1388), .Z(n1386) );
  NAND U1617 ( .A(n556), .B(msg[15]), .Z(n1388) );
  AND U1618 ( .A(n1389), .B(n1390), .Z(n1387) );
  NAND U1619 ( .A(n1391), .B(n560), .Z(n1390) );
  XOR U1620 ( .A(n1392), .B(n1393), .Z(n1391) );
  XOR U1621 ( .A(n2615), .B(n1276), .Z(n1393) );
  IV U1622 ( .A(n1304), .Z(n1276) );
  XNOR U1623 ( .A(shift_row_out[31]), .B(shift_row_out[7]), .Z(n1304) );
  XNOR U1624 ( .A(shift_row_out[23]), .B(n779), .Z(n1392) );
  IV U1625 ( .A(n2210), .Z(n779) );
  NAND U1626 ( .A(shift_row_out[15]), .B(n566), .Z(n1389) );
  XOR U1627 ( .A(n1394), .B(key[14]), .Z(o[14]) );
  NAND U1628 ( .A(n1395), .B(n1396), .Z(n1394) );
  NAND U1629 ( .A(n556), .B(msg[14]), .Z(n1396) );
  AND U1630 ( .A(n1397), .B(n1398), .Z(n1395) );
  NAND U1631 ( .A(n1399), .B(n560), .Z(n1398) );
  XOR U1632 ( .A(n1400), .B(n1401), .Z(n1399) );
  XNOR U1633 ( .A(n1265), .B(n2615), .Z(n1401) );
  IV U1634 ( .A(n2209), .Z(n1265) );
  XOR U1635 ( .A(n2614), .B(n1238), .Z(n1400) );
  NANDN U1636 ( .B(n2210), .A(n566), .Z(n1397) );
  XOR U1637 ( .A(n1402), .B(key[13]), .Z(o[13]) );
  NAND U1638 ( .A(n1403), .B(n1404), .Z(n1402) );
  NAND U1639 ( .A(n556), .B(msg[13]), .Z(n1404) );
  AND U1640 ( .A(n1405), .B(n1406), .Z(n1403) );
  NAND U1641 ( .A(n1407), .B(n560), .Z(n1406) );
  XOR U1642 ( .A(n1408), .B(n1409), .Z(n1407) );
  XOR U1643 ( .A(shift_row_out[20]), .B(shift_row_out[12]), .Z(n1409) );
  XOR U1644 ( .A(n2614), .B(n1247), .Z(n1408) );
  XNOR U1645 ( .A(\b/SBOX[0].sbox/n90 ), .B(n3019), .Z(n1247) );
  NANDN U1646 ( .B(n2209), .A(n566), .Z(n1405) );
  XOR U1647 ( .A(n1410), .B(key[12]), .Z(o[12]) );
  NAND U1648 ( .A(n1411), .B(n1412), .Z(n1410) );
  NAND U1649 ( .A(n556), .B(msg[12]), .Z(n1412) );
  AND U1650 ( .A(n1413), .B(n1414), .Z(n1411) );
  NAND U1651 ( .A(n1415), .B(n560), .Z(n1414) );
  XOR U1652 ( .A(n1416), .B(n1417), .Z(n1415) );
  XNOR U1653 ( .A(n564), .B(n1266), .Z(n1417) );
  XNOR U1654 ( .A(shift_row_out[28]), .B(shift_row_out[4]), .Z(n1266) );
  XOR U1655 ( .A(shift_row_out[11]), .B(n1418), .Z(n1416) );
  XOR U1656 ( .A(shift_row_out[20]), .B(shift_row_out[19]), .Z(n1418) );
  NAND U1657 ( .A(n566), .B(shift_row_out[12]), .Z(n1413) );
  XOR U1658 ( .A(n1419), .B(key[127]), .Z(o[127]) );
  NAND U1659 ( .A(n1420), .B(n1421), .Z(n1419) );
  NAND U1660 ( .A(n556), .B(msg[127]), .Z(n1421) );
  AND U1661 ( .A(n1422), .B(n1423), .Z(n1420) );
  NAND U1662 ( .A(n1424), .B(n560), .Z(n1423) );
  XOR U1663 ( .A(n1425), .B(n1426), .Z(n1424) );
  XOR U1664 ( .A(n2696), .B(n1427), .Z(n1426) );
  XNOR U1665 ( .A(shift_row_out[103]), .B(n1428), .Z(n1425) );
  NAND U1666 ( .A(n566), .B(shift_row_out[127]), .Z(n1422) );
  XOR U1667 ( .A(n1429), .B(key[126]), .Z(o[126]) );
  NAND U1668 ( .A(n1430), .B(n1431), .Z(n1429) );
  NAND U1669 ( .A(n556), .B(msg[126]), .Z(n1431) );
  AND U1670 ( .A(n1432), .B(n1433), .Z(n1430) );
  NAND U1671 ( .A(n1434), .B(n560), .Z(n1433) );
  XOR U1672 ( .A(n1435), .B(n1436), .Z(n1434) );
  XNOR U1673 ( .A(n1428), .B(n2776), .Z(n1436) );
  XOR U1674 ( .A(n2695), .B(n1437), .Z(n1435) );
  NANDN U1675 ( .B(n2696), .A(n566), .Z(n1432) );
  XOR U1676 ( .A(n1438), .B(key[125]), .Z(o[125]) );
  NAND U1677 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U1678 ( .A(n556), .B(msg[125]), .Z(n1440) );
  AND U1679 ( .A(n1441), .B(n1442), .Z(n1439) );
  NAND U1680 ( .A(n1443), .B(n560), .Z(n1442) );
  XOR U1681 ( .A(n1444), .B(n1445), .Z(n1443) );
  XOR U1682 ( .A(shift_row_out[124]), .B(shift_row_out[100]), .Z(n1445) );
  XOR U1683 ( .A(n2776), .B(n1446), .Z(n1444) );
  NANDN U1684 ( .B(n2695), .A(n566), .Z(n1441) );
  XOR U1685 ( .A(n1447), .B(key[124]), .Z(o[124]) );
  NAND U1686 ( .A(n1448), .B(n1449), .Z(n1447) );
  NAND U1687 ( .A(n556), .B(msg[124]), .Z(n1449) );
  AND U1688 ( .A(n1450), .B(n1451), .Z(n1448) );
  NAND U1689 ( .A(n1452), .B(n560), .Z(n1451) );
  XOR U1690 ( .A(n1453), .B(n1454), .Z(n1452) );
  XOR U1691 ( .A(n1455), .B(n1456), .Z(n1454) );
  XNOR U1692 ( .A(shift_row_out[100]), .B(n1457), .Z(n1453) );
  NAND U1693 ( .A(n566), .B(shift_row_out[124]), .Z(n1450) );
  XOR U1694 ( .A(n1458), .B(key[123]), .Z(o[123]) );
  NAND U1695 ( .A(n1459), .B(n1460), .Z(n1458) );
  NAND U1696 ( .A(n556), .B(msg[123]), .Z(n1460) );
  AND U1697 ( .A(n1461), .B(n1462), .Z(n1459) );
  NAND U1698 ( .A(n1463), .B(n560), .Z(n1462) );
  XOR U1699 ( .A(n1464), .B(n1465), .Z(n1463) );
  XOR U1700 ( .A(n1455), .B(n1466), .Z(n1465) );
  XOR U1701 ( .A(shift_row_out[107]), .B(n1467), .Z(n1464) );
  XOR U1702 ( .A(shift_row_out[99]), .B(shift_row_out[115]), .Z(n1467) );
  NAND U1703 ( .A(n566), .B(shift_row_out[123]), .Z(n1461) );
  XOR U1704 ( .A(n1468), .B(key[122]), .Z(o[122]) );
  NAND U1705 ( .A(n1469), .B(n1470), .Z(n1468) );
  NAND U1706 ( .A(msg[122]), .B(n556), .Z(n1470) );
  AND U1707 ( .A(n1471), .B(n1472), .Z(n1469) );
  NAND U1708 ( .A(n1473), .B(n560), .Z(n1472) );
  XOR U1709 ( .A(n1474), .B(n1475), .Z(n1473) );
  XNOR U1710 ( .A(shift_row_out[106]), .B(n1476), .Z(n1475) );
  XOR U1711 ( .A(shift_row_out[98]), .B(shift_row_out[114]), .Z(n1474) );
  NAND U1712 ( .A(n566), .B(shift_row_out[122]), .Z(n1471) );
  XOR U1713 ( .A(n1477), .B(key[121]), .Z(o[121]) );
  NAND U1714 ( .A(n1478), .B(n1479), .Z(n1477) );
  NAND U1715 ( .A(n556), .B(msg[121]), .Z(n1479) );
  AND U1716 ( .A(n1480), .B(n1481), .Z(n1478) );
  NAND U1717 ( .A(n1482), .B(n560), .Z(n1481) );
  XOR U1718 ( .A(n1483), .B(n1484), .Z(n1482) );
  XNOR U1719 ( .A(n1455), .B(n1485), .Z(n1484) );
  XNOR U1720 ( .A(n2775), .B(n1486), .Z(n1483) );
  XNOR U1721 ( .A(n2289), .B(n587), .Z(n1486) );
  NANDN U1722 ( .B(n2694), .A(n566), .Z(n1480) );
  XOR U1723 ( .A(n1487), .B(key[120]), .Z(o[120]) );
  NAND U1724 ( .A(n1488), .B(n1489), .Z(n1487) );
  NAND U1725 ( .A(n556), .B(msg[120]), .Z(n1489) );
  AND U1726 ( .A(n1490), .B(n1491), .Z(n1488) );
  NAND U1727 ( .A(n1492), .B(n560), .Z(n1491) );
  XOR U1728 ( .A(n1493), .B(n1494), .Z(n1492) );
  XNOR U1729 ( .A(n1495), .B(n1883), .Z(n1494) );
  XOR U1730 ( .A(n2774), .B(n1455), .Z(n1493) );
  XNOR U1731 ( .A(shift_row_out[103]), .B(shift_row_out[127]), .Z(n1455) );
  NANDN U1732 ( .B(n2693), .A(n566), .Z(n1490) );
  XOR U1733 ( .A(n1496), .B(key[11]), .Z(o[11]) );
  NAND U1734 ( .A(n1497), .B(n1498), .Z(n1496) );
  NAND U1735 ( .A(n556), .B(msg[11]), .Z(n1498) );
  AND U1736 ( .A(n1499), .B(n1500), .Z(n1497) );
  NAND U1737 ( .A(n1501), .B(n560), .Z(n1500) );
  XOR U1738 ( .A(n1502), .B(n1503), .Z(n1501) );
  XNOR U1739 ( .A(n564), .B(n1275), .Z(n1503) );
  XNOR U1740 ( .A(shift_row_out[27]), .B(shift_row_out[3]), .Z(n1275) );
  XOR U1741 ( .A(shift_row_out[15]), .B(shift_row_out[23]), .Z(n564) );
  XOR U1742 ( .A(shift_row_out[10]), .B(n1504), .Z(n1502) );
  XOR U1743 ( .A(shift_row_out[19]), .B(shift_row_out[18]), .Z(n1504) );
  NAND U1744 ( .A(n566), .B(shift_row_out[11]), .Z(n1499) );
  XOR U1745 ( .A(n1505), .B(key[119]), .Z(o[119]) );
  NAND U1746 ( .A(n1506), .B(n1507), .Z(n1505) );
  NAND U1747 ( .A(n556), .B(msg[119]), .Z(n1507) );
  AND U1748 ( .A(n1508), .B(n1509), .Z(n1506) );
  NAND U1749 ( .A(n1510), .B(n560), .Z(n1509) );
  XOR U1750 ( .A(n1511), .B(n1512), .Z(n1510) );
  XNOR U1751 ( .A(shift_row_out[103]), .B(n1513), .Z(n1512) );
  XOR U1752 ( .A(shift_row_out[127]), .B(shift_row_out[111]), .Z(n1511) );
  NAND U1753 ( .A(n566), .B(shift_row_out[119]), .Z(n1508) );
  XOR U1754 ( .A(n1514), .B(key[118]), .Z(o[118]) );
  NAND U1755 ( .A(n1515), .B(n1516), .Z(n1514) );
  NAND U1756 ( .A(n556), .B(msg[118]), .Z(n1516) );
  AND U1757 ( .A(n1517), .B(n1518), .Z(n1515) );
  NAND U1758 ( .A(n1519), .B(n560), .Z(n1518) );
  XOR U1759 ( .A(n1520), .B(n1521), .Z(n1519) );
  XNOR U1760 ( .A(n1522), .B(n2777), .Z(n1521) );
  XOR U1761 ( .A(n2696), .B(n1523), .Z(n1520) );
  NANDN U1762 ( .B(n2291), .A(n566), .Z(n1517) );
  XOR U1763 ( .A(n1524), .B(key[117]), .Z(o[117]) );
  NAND U1764 ( .A(n1525), .B(n1526), .Z(n1524) );
  NAND U1765 ( .A(n556), .B(msg[117]), .Z(n1526) );
  AND U1766 ( .A(n1527), .B(n1528), .Z(n1525) );
  NAND U1767 ( .A(n1529), .B(n560), .Z(n1528) );
  XOR U1768 ( .A(n1530), .B(n1531), .Z(n1529) );
  XOR U1769 ( .A(n2695), .B(n1532), .Z(n1530) );
  NANDN U1770 ( .B(n2290), .A(n566), .Z(n1527) );
  XOR U1771 ( .A(n1533), .B(key[116]), .Z(o[116]) );
  NAND U1772 ( .A(n1534), .B(n1535), .Z(n1533) );
  NAND U1773 ( .A(n556), .B(msg[116]), .Z(n1535) );
  AND U1774 ( .A(n1536), .B(n1537), .Z(n1534) );
  NAND U1775 ( .A(n1538), .B(n560), .Z(n1537) );
  XOR U1776 ( .A(n1539), .B(n1540), .Z(n1538) );
  XOR U1777 ( .A(n576), .B(n1541), .Z(n1540) );
  XNOR U1778 ( .A(shift_row_out[115]), .B(shift_row_out[123]), .Z(n576) );
  XOR U1779 ( .A(shift_row_out[100]), .B(n1542), .Z(n1539) );
  XOR U1780 ( .A(shift_row_out[124]), .B(shift_row_out[108]), .Z(n1542) );
  NAND U1781 ( .A(n566), .B(shift_row_out[116]), .Z(n1536) );
  XOR U1782 ( .A(n1543), .B(key[115]), .Z(o[115]) );
  NAND U1783 ( .A(n1544), .B(n1545), .Z(n1543) );
  NAND U1784 ( .A(n556), .B(msg[115]), .Z(n1545) );
  AND U1785 ( .A(n1546), .B(n1547), .Z(n1544) );
  NAND U1786 ( .A(n1548), .B(n560), .Z(n1547) );
  XOR U1787 ( .A(n1549), .B(n1550), .Z(n1548) );
  XOR U1788 ( .A(n1457), .B(n1541), .Z(n1550) );
  XNOR U1789 ( .A(shift_row_out[107]), .B(n586), .Z(n1549) );
  XNOR U1790 ( .A(shift_row_out[114]), .B(shift_row_out[122]), .Z(n586) );
  NAND U1791 ( .A(n566), .B(shift_row_out[115]), .Z(n1546) );
  XOR U1792 ( .A(n1551), .B(key[114]), .Z(o[114]) );
  NAND U1793 ( .A(n1552), .B(n1553), .Z(n1551) );
  NAND U1794 ( .A(msg[114]), .B(n556), .Z(n1553) );
  AND U1795 ( .A(n1554), .B(n1555), .Z(n1552) );
  NAND U1796 ( .A(n1556), .B(n560), .Z(n1555) );
  XNOR U1797 ( .A(n1466), .B(n1557), .Z(n1556) );
  XNOR U1798 ( .A(shift_row_out[106]), .B(n596), .Z(n1557) );
  XNOR U1799 ( .A(n2694), .B(n2289), .Z(n596) );
  NAND U1800 ( .A(n566), .B(shift_row_out[114]), .Z(n1554) );
  XOR U1801 ( .A(n1558), .B(key[113]), .Z(o[113]) );
  NAND U1802 ( .A(n1559), .B(n1560), .Z(n1558) );
  NAND U1803 ( .A(n556), .B(msg[113]), .Z(n1560) );
  AND U1804 ( .A(n1561), .B(n1562), .Z(n1559) );
  NAND U1805 ( .A(n1563), .B(n560), .Z(n1562) );
  XOR U1806 ( .A(n1564), .B(n1565), .Z(n1563) );
  XOR U1807 ( .A(n1476), .B(n1541), .Z(n1565) );
  XOR U1808 ( .A(n1884), .B(n605), .Z(n1564) );
  XNOR U1809 ( .A(n2693), .B(n2288), .Z(n605) );
  NANDN U1810 ( .B(n2289), .A(n566), .Z(n1561) );
  XOR U1811 ( .A(n1566), .B(key[112]), .Z(o[112]) );
  NAND U1812 ( .A(n1567), .B(n1568), .Z(n1566) );
  NAND U1813 ( .A(n556), .B(msg[112]), .Z(n1568) );
  AND U1814 ( .A(n1569), .B(n1570), .Z(n1567) );
  NAND U1815 ( .A(n1571), .B(n560), .Z(n1570) );
  XNOR U1816 ( .A(n1572), .B(n1541), .Z(n1571) );
  XNOR U1817 ( .A(n1883), .B(n1485), .Z(n1572) );
  NANDN U1818 ( .B(n2288), .A(n566), .Z(n1569) );
  XOR U1819 ( .A(n1573), .B(key[111]), .Z(o[111]) );
  NAND U1820 ( .A(n1574), .B(n1575), .Z(n1573) );
  NAND U1821 ( .A(n556), .B(msg[111]), .Z(n1575) );
  AND U1822 ( .A(n1576), .B(n1577), .Z(n1574) );
  NAND U1823 ( .A(n1578), .B(n560), .Z(n1577) );
  XNOR U1824 ( .A(n1541), .B(n1579), .Z(n1578) );
  XNOR U1825 ( .A(shift_row_out[103]), .B(n1437), .Z(n1579) );
  XNOR U1826 ( .A(n1886), .B(n2291), .Z(n1437) );
  NAND U1827 ( .A(n566), .B(shift_row_out[111]), .Z(n1576) );
  XOR U1828 ( .A(n1580), .B(key[110]), .Z(o[110]) );
  NAND U1829 ( .A(n1581), .B(n1582), .Z(n1580) );
  NAND U1830 ( .A(n556), .B(msg[110]), .Z(n1582) );
  AND U1831 ( .A(n1583), .B(n1584), .Z(n1581) );
  NAND U1832 ( .A(n1585), .B(n560), .Z(n1584) );
  XNOR U1833 ( .A(n1586), .B(n1513), .Z(n1585) );
  XOR U1834 ( .A(n2777), .B(n1446), .Z(n1586) );
  XNOR U1835 ( .A(n1885), .B(n2290), .Z(n1446) );
  NANDN U1836 ( .B(n1886), .A(n566), .Z(n1583) );
  XOR U1837 ( .A(n1587), .B(key[10]), .Z(o[10]) );
  NAND U1838 ( .A(n1588), .B(n1589), .Z(n1587) );
  NAND U1839 ( .A(msg[10]), .B(n556), .Z(n1589) );
  AND U1840 ( .A(n1590), .B(n1591), .Z(n1588) );
  NAND U1841 ( .A(n1592), .B(n560), .Z(n1591) );
  XOR U1842 ( .A(n1593), .B(n1369), .Z(n1592) );
  XOR U1843 ( .A(n1353), .B(n1286), .Z(n1369) );
  XNOR U1844 ( .A(shift_row_out[26]), .B(shift_row_out[2]), .Z(n1286) );
  IV U1845 ( .A(n2613), .Z(n1353) );
  XOR U1846 ( .A(shift_row_out[18]), .B(n2208), .Z(n1593) );
  NAND U1847 ( .A(n566), .B(shift_row_out[10]), .Z(n1590) );
  XOR U1848 ( .A(n1594), .B(key[109]), .Z(o[109]) );
  NAND U1849 ( .A(n1595), .B(n1596), .Z(n1594) );
  NAND U1850 ( .A(n556), .B(msg[109]), .Z(n1596) );
  AND U1851 ( .A(n1597), .B(n1598), .Z(n1595) );
  NAND U1852 ( .A(n1599), .B(n560), .Z(n1598) );
  XNOR U1853 ( .A(n1600), .B(n1523), .Z(n1599) );
  XOR U1854 ( .A(n2776), .B(n1456), .Z(n1600) );
  XNOR U1855 ( .A(shift_row_out[108]), .B(shift_row_out[116]), .Z(n1456) );
  NANDN U1856 ( .B(n1885), .A(n566), .Z(n1597) );
  XOR U1857 ( .A(n1601), .B(key[108]), .Z(o[108]) );
  NAND U1858 ( .A(n1602), .B(n1603), .Z(n1601) );
  NAND U1859 ( .A(n556), .B(msg[108]), .Z(n1603) );
  AND U1860 ( .A(n1604), .B(n1605), .Z(n1602) );
  NAND U1861 ( .A(n1606), .B(n560), .Z(n1605) );
  XOR U1862 ( .A(n1607), .B(n1608), .Z(n1606) );
  XOR U1863 ( .A(n1609), .B(n1532), .Z(n1608) );
  XOR U1864 ( .A(shift_row_out[100]), .B(n1610), .Z(n1607) );
  XOR U1865 ( .A(shift_row_out[115]), .B(shift_row_out[107]), .Z(n1610) );
  NAND U1866 ( .A(n566), .B(shift_row_out[108]), .Z(n1604) );
  XOR U1867 ( .A(n1611), .B(key[107]), .Z(o[107]) );
  NAND U1868 ( .A(n1612), .B(n1613), .Z(n1611) );
  NAND U1869 ( .A(n556), .B(msg[107]), .Z(n1613) );
  AND U1870 ( .A(n1614), .B(n1615), .Z(n1612) );
  NAND U1871 ( .A(n1616), .B(n560), .Z(n1615) );
  XOR U1872 ( .A(n1617), .B(n1618), .Z(n1616) );
  XOR U1873 ( .A(n1609), .B(n1457), .Z(n1618) );
  XNOR U1874 ( .A(shift_row_out[123]), .B(shift_row_out[99]), .Z(n1457) );
  XOR U1875 ( .A(shift_row_out[106]), .B(n1619), .Z(n1617) );
  XOR U1876 ( .A(shift_row_out[115]), .B(shift_row_out[114]), .Z(n1619) );
  NAND U1877 ( .A(n566), .B(shift_row_out[107]), .Z(n1614) );
  XOR U1878 ( .A(n1620), .B(key[106]), .Z(o[106]) );
  NAND U1879 ( .A(n1621), .B(n1622), .Z(n1620) );
  NAND U1880 ( .A(msg[106]), .B(n556), .Z(n1622) );
  AND U1881 ( .A(n1623), .B(n1624), .Z(n1621) );
  NAND U1882 ( .A(n1625), .B(n560), .Z(n1624) );
  XOR U1883 ( .A(n1626), .B(n1627), .Z(n1625) );
  XOR U1884 ( .A(n587), .B(n1466), .Z(n1627) );
  XNOR U1885 ( .A(shift_row_out[122]), .B(shift_row_out[98]), .Z(n1466) );
  IV U1886 ( .A(n1884), .Z(n587) );
  XOR U1887 ( .A(shift_row_out[114]), .B(n2289), .Z(n1626) );
  NAND U1888 ( .A(n566), .B(shift_row_out[106]), .Z(n1623) );
  XOR U1889 ( .A(n1628), .B(key[105]), .Z(o[105]) );
  NAND U1890 ( .A(n1629), .B(n1630), .Z(n1628) );
  NAND U1891 ( .A(n556), .B(msg[105]), .Z(n1630) );
  AND U1892 ( .A(n1631), .B(n1632), .Z(n1629) );
  NAND U1893 ( .A(n1633), .B(n560), .Z(n1632) );
  XOR U1894 ( .A(n1634), .B(n1635), .Z(n1633) );
  XNOR U1895 ( .A(n1427), .B(n1476), .Z(n1635) );
  XNOR U1896 ( .A(n1883), .B(n1636), .Z(n1634) );
  XNOR U1897 ( .A(n2289), .B(n1495), .Z(n1636) );
  IV U1898 ( .A(n2288), .Z(n1495) );
  NANDN U1899 ( .B(n1884), .A(n566), .Z(n1631) );
  XOR U1900 ( .A(n1637), .B(key[104]), .Z(o[104]) );
  NAND U1901 ( .A(n1638), .B(n1639), .Z(n1637) );
  NAND U1902 ( .A(n556), .B(msg[104]), .Z(n1639) );
  AND U1903 ( .A(n1640), .B(n1641), .Z(n1638) );
  NAND U1904 ( .A(n1642), .B(n560), .Z(n1641) );
  XOR U1905 ( .A(n1643), .B(n1485), .Z(n1642) );
  XOR U1906 ( .A(n2288), .B(n1609), .Z(n1643) );
  IV U1907 ( .A(n1427), .Z(n1609) );
  XOR U1908 ( .A(shift_row_out[111]), .B(shift_row_out[119]), .Z(n1427) );
  NANDN U1909 ( .B(n1883), .A(n566), .Z(n1640) );
  XOR U1910 ( .A(n1644), .B(key[103]), .Z(o[103]) );
  NAND U1911 ( .A(n1645), .B(n1646), .Z(n1644) );
  NAND U1912 ( .A(msg[103]), .B(n556), .Z(n1646) );
  AND U1913 ( .A(n1647), .B(n1648), .Z(n1645) );
  NAND U1914 ( .A(n1649), .B(n560), .Z(n1648) );
  XOR U1915 ( .A(n1650), .B(n1651), .Z(n1649) );
  XOR U1916 ( .A(n1428), .B(n1541), .Z(n1651) );
  XNOR U1917 ( .A(shift_row_out[119]), .B(shift_row_out[127]), .Z(n1541) );
  IV U1918 ( .A(n2777), .Z(n1428) );
  XNOR U1919 ( .A(shift_row_out[111]), .B(n1522), .Z(n1650) );
  NAND U1920 ( .A(n566), .B(shift_row_out[103]), .Z(n1647) );
  XOR U1921 ( .A(n1652), .B(key[102]), .Z(o[102]) );
  NAND U1922 ( .A(n1653), .B(n1654), .Z(n1652) );
  NAND U1923 ( .A(n556), .B(msg[102]), .Z(n1654) );
  AND U1924 ( .A(n1655), .B(n1656), .Z(n1653) );
  NAND U1925 ( .A(n1657), .B(n560), .Z(n1656) );
  XOR U1926 ( .A(n1658), .B(n1659), .Z(n1657) );
  XNOR U1927 ( .A(n1522), .B(n1885), .Z(n1659) );
  IV U1928 ( .A(n1886), .Z(n1522) );
  XOR U1929 ( .A(n2776), .B(n1513), .Z(n1658) );
  NANDN U1930 ( .B(n2777), .A(n566), .Z(n1655) );
  XOR U1931 ( .A(n1660), .B(key[101]), .Z(o[101]) );
  NAND U1932 ( .A(n1661), .B(n1662), .Z(n1660) );
  NAND U1933 ( .A(n556), .B(msg[101]), .Z(n1662) );
  AND U1934 ( .A(n1663), .B(n1664), .Z(n1661) );
  NAND U1935 ( .A(n1665), .B(n560), .Z(n1664) );
  XOR U1936 ( .A(n1666), .B(n1667), .Z(n1665) );
  XOR U1937 ( .A(shift_row_out[108]), .B(shift_row_out[100]), .Z(n1667) );
  XOR U1938 ( .A(n1885), .B(n1523), .Z(n1666) );
  XNOR U1939 ( .A(n2695), .B(n2290), .Z(n1523) );
  NANDN U1940 ( .B(n2776), .A(n566), .Z(n1663) );
  XOR U1941 ( .A(n1668), .B(key[100]), .Z(o[100]) );
  NAND U1942 ( .A(n1669), .B(n1670), .Z(n1668) );
  NAND U1943 ( .A(msg[100]), .B(n556), .Z(n1670) );
  AND U1944 ( .A(n1671), .B(n1672), .Z(n1669) );
  NAND U1945 ( .A(n1673), .B(n560), .Z(n1672) );
  XOR U1946 ( .A(n1674), .B(n1675), .Z(n1673) );
  XNOR U1947 ( .A(n606), .B(n1532), .Z(n1675) );
  XNOR U1948 ( .A(shift_row_out[116]), .B(shift_row_out[124]), .Z(n1532) );
  XOR U1949 ( .A(shift_row_out[103]), .B(shift_row_out[111]), .Z(n606) );
  XOR U1950 ( .A(shift_row_out[107]), .B(n1676), .Z(n1674) );
  XOR U1951 ( .A(shift_row_out[99]), .B(shift_row_out[108]), .Z(n1676) );
  NAND U1952 ( .A(n566), .B(shift_row_out[100]), .Z(n1671) );
  XOR U1953 ( .A(n1677), .B(key[0]), .Z(o[0]) );
  NAND U1954 ( .A(n1678), .B(n1679), .Z(n1677) );
  NAND U1955 ( .A(msg[0]), .B(n556), .Z(n1679) );
  AND U1956 ( .A(n1680), .B(n1681), .Z(n1678) );
  NAND U1957 ( .A(n1682), .B(n560), .Z(n1681) );
  NOR U1958 ( .A(n556), .B(n566), .Z(n560) );
  AND U1959 ( .A(n1683), .B(n1684), .Z(n556) );
  ANDN U1960 ( .A(n1685), .B(counter[3]), .Z(n1684) );
  XNOR U1961 ( .A(n1686), .B(n1385), .Z(n1682) );
  XNOR U1962 ( .A(n3017), .B(n2207), .Z(n1385) );
  XOR U1963 ( .A(n2612), .B(n1070), .Z(n1686) );
  XNOR U1964 ( .A(shift_row_out[15]), .B(shift_row_out[7]), .Z(n1070) );
  NANDN U1965 ( .B(\b/SBOX[0].sbox/n88 ), .A(n566), .Z(n1680) );
  XNOR U1966 ( .A(\e/n97 ), .B(n539), .Z(nextKey[9]) );
  IV U1967 ( .A(\e/n291 ), .Z(nextKey[95]) );
  IV U1968 ( .A(\e/n290 ), .Z(nextKey[94]) );
  IV U1969 ( .A(\e/n289 ), .Z(nextKey[93]) );
  IV U1970 ( .A(\e/n288 ), .Z(nextKey[92]) );
  IV U1971 ( .A(\e/n287 ), .Z(nextKey[91]) );
  IV U1972 ( .A(\e/n286 ), .Z(nextKey[90]) );
  XNOR U1973 ( .A(\e/n98 ), .B(n540), .Z(nextKey[8]) );
  IV U1974 ( .A(\e/n285 ), .Z(nextKey[89]) );
  IV U1975 ( .A(\e/n284 ), .Z(nextKey[88]) );
  IV U1976 ( .A(\e/n283 ), .Z(nextKey[87]) );
  IV U1977 ( .A(\e/n282 ), .Z(nextKey[86]) );
  IV U1978 ( .A(\e/n281 ), .Z(nextKey[85]) );
  IV U1979 ( .A(\e/n280 ), .Z(nextKey[84]) );
  IV U1980 ( .A(\e/n279 ), .Z(nextKey[83]) );
  IV U1981 ( .A(\e/n278 ), .Z(nextKey[82]) );
  IV U1982 ( .A(\e/n277 ), .Z(nextKey[81]) );
  IV U1983 ( .A(\e/n276 ), .Z(nextKey[80]) );
  IV U1984 ( .A(\e/n275 ), .Z(nextKey[79]) );
  IV U1985 ( .A(\e/n274 ), .Z(nextKey[78]) );
  IV U1986 ( .A(\e/n273 ), .Z(nextKey[77]) );
  IV U1987 ( .A(\e/n272 ), .Z(nextKey[76]) );
  IV U1988 ( .A(\e/n271 ), .Z(nextKey[75]) );
  IV U1989 ( .A(\e/n270 ), .Z(nextKey[74]) );
  IV U1990 ( .A(\e/n269 ), .Z(nextKey[73]) );
  IV U1991 ( .A(\e/n268 ), .Z(nextKey[72]) );
  IV U1992 ( .A(\e/n267 ), .Z(nextKey[39]) );
  IV U1993 ( .A(\e/n266 ), .Z(nextKey[38]) );
  IV U1994 ( .A(\e/n265 ), .Z(nextKey[37]) );
  IV U1995 ( .A(\e/n264 ), .Z(nextKey[36]) );
  IV U1996 ( .A(\e/n263 ), .Z(nextKey[35]) );
  IV U1997 ( .A(\e/n262 ), .Z(nextKey[34]) );
  IV U1998 ( .A(\e/n261 ), .Z(nextKey[33]) );
  IV U1999 ( .A(\e/n260 ), .Z(nextKey[32]) );
  XNOR U2000 ( .A(\e/t[31] ), .B(\e/n75 ), .Z(nextKey[31]) );
  XNOR U2001 ( .A(\e/n76 ), .B(n529), .Z(nextKey[30]) );
  XNOR U2002 ( .A(\e/n77 ), .B(n530), .Z(nextKey[29]) );
  XNOR U2003 ( .A(\e/t[28] ), .B(\e/n78 ), .Z(nextKey[28]) );
  XNOR U2004 ( .A(\e/t[27] ), .B(\e/n79 ), .Z(nextKey[27]) );
  XNOR U2005 ( .A(\e/t[26] ), .B(\e/n80 ), .Z(nextKey[26]) );
  XNOR U2006 ( .A(\e/n81 ), .B(n531), .Z(nextKey[25]) );
  XNOR U2007 ( .A(\e/n82 ), .B(n532), .Z(nextKey[24]) );
  XNOR U2008 ( .A(\e/t[23] ), .B(\e/n83 ), .Z(nextKey[23]) );
  XNOR U2009 ( .A(\e/n84 ), .B(n533), .Z(nextKey[22]) );
  XNOR U2010 ( .A(\e/n85 ), .B(n534), .Z(nextKey[21]) );
  XNOR U2011 ( .A(\e/t[20] ), .B(\e/n86 ), .Z(nextKey[20]) );
  XNOR U2012 ( .A(\e/t[19] ), .B(\e/n87 ), .Z(nextKey[19]) );
  XNOR U2013 ( .A(\e/t[18] ), .B(\e/n88 ), .Z(nextKey[18]) );
  XNOR U2014 ( .A(\e/n89 ), .B(n535), .Z(nextKey[17]) );
  XNOR U2015 ( .A(\e/n90 ), .B(n536), .Z(nextKey[16]) );
  XNOR U2016 ( .A(\e/t[15] ), .B(\e/n91 ), .Z(nextKey[15]) );
  XNOR U2017 ( .A(\e/n92 ), .B(n537), .Z(nextKey[14]) );
  XNOR U2018 ( .A(\e/n93 ), .B(n538), .Z(nextKey[13]) );
  XNOR U2019 ( .A(\e/t[12] ), .B(\e/n94 ), .Z(nextKey[12]) );
  XNOR U2020 ( .A(\e/t[11] ), .B(\e/n95 ), .Z(nextKey[11]) );
  XNOR U2021 ( .A(\e/t[10] ), .B(\e/n96 ), .Z(nextKey[10]) );
  NANDN U2022 ( .B(n566), .A(key[8]), .Z(\e/n98 ) );
  NANDN U2023 ( .B(n566), .A(key[9]), .Z(\e/n97 ) );
  NANDN U2024 ( .B(n566), .A(key[10]), .Z(\e/n96 ) );
  NANDN U2025 ( .B(n566), .A(key[11]), .Z(\e/n95 ) );
  NANDN U2026 ( .B(n566), .A(key[12]), .Z(\e/n94 ) );
  NANDN U2027 ( .B(n566), .A(key[13]), .Z(\e/n93 ) );
  NANDN U2028 ( .B(n566), .A(key[14]), .Z(\e/n92 ) );
  NANDN U2029 ( .B(n566), .A(key[15]), .Z(\e/n91 ) );
  NANDN U2030 ( .B(n566), .A(key[16]), .Z(\e/n90 ) );
  NANDN U2031 ( .B(n566), .A(key[17]), .Z(\e/n89 ) );
  NANDN U2032 ( .B(n566), .A(key[18]), .Z(\e/n88 ) );
  NANDN U2033 ( .B(n566), .A(key[19]), .Z(\e/n87 ) );
  NANDN U2034 ( .B(n566), .A(key[20]), .Z(\e/n86 ) );
  NANDN U2035 ( .B(n566), .A(key[21]), .Z(\e/n85 ) );
  NANDN U2036 ( .B(n566), .A(key[22]), .Z(\e/n84 ) );
  NANDN U2037 ( .B(n566), .A(key[23]), .Z(\e/n83 ) );
  NANDN U2038 ( .B(n566), .A(key[24]), .Z(\e/n82 ) );
  NANDN U2039 ( .B(n566), .A(key[25]), .Z(\e/n81 ) );
  NANDN U2040 ( .B(n566), .A(key[26]), .Z(\e/n80 ) );
  NANDN U2041 ( .B(n566), .A(key[27]), .Z(\e/n79 ) );
  NANDN U2042 ( .B(n566), .A(key[28]), .Z(\e/n78 ) );
  NANDN U2043 ( .B(n566), .A(key[29]), .Z(\e/n77 ) );
  NANDN U2044 ( .B(n566), .A(key[30]), .Z(\e/n76 ) );
  NANDN U2045 ( .B(n566), .A(key[31]), .Z(\e/n75 ) );
  AND U2046 ( .A(key[99]), .B(n1687), .Z(\e/w[3][3] ) );
  AND U2047 ( .A(key[101]), .B(n1687), .Z(\e/w[3][5] ) );
  AND U2048 ( .A(key[102]), .B(n1687), .Z(\e/w[3][6] ) );
  AND U2049 ( .A(key[107]), .B(n1687), .Z(\e/w[3][11] ) );
  AND U2050 ( .A(key[109]), .B(n1687), .Z(\e/w[3][13] ) );
  AND U2051 ( .A(key[110]), .B(n1687), .Z(\e/w[3][14] ) );
  AND U2052 ( .A(key[115]), .B(n1687), .Z(\e/w[3][19] ) );
  AND U2053 ( .A(key[117]), .B(n1687), .Z(\e/w[3][21] ) );
  AND U2054 ( .A(key[118]), .B(n1687), .Z(\e/w[3][22] ) );
  AND U2055 ( .A(key[123]), .B(n1687), .Z(\e/w[3][27] ) );
  AND U2056 ( .A(key[125]), .B(n1687), .Z(\e/w[3][29] ) );
  AND U2057 ( .A(key[126]), .B(n1687), .Z(\e/w[3][30] ) );
  NANDN U2058 ( .B(n566), .A(key[95]), .Z(\e/n259 ) );
  NANDN U2059 ( .B(n566), .A(key[94]), .Z(\e/n258 ) );
  NANDN U2060 ( .B(n566), .A(key[93]), .Z(\e/n257 ) );
  NANDN U2061 ( .B(n566), .A(key[92]), .Z(\e/n256 ) );
  NANDN U2062 ( .B(n566), .A(key[91]), .Z(\e/n255 ) );
  NANDN U2063 ( .B(n566), .A(key[90]), .Z(\e/n254 ) );
  NANDN U2064 ( .B(n566), .A(key[89]), .Z(\e/n253 ) );
  NANDN U2065 ( .B(n566), .A(key[88]), .Z(\e/n252 ) );
  NANDN U2066 ( .B(n566), .A(key[87]), .Z(\e/n251 ) );
  NANDN U2067 ( .B(n566), .A(key[86]), .Z(\e/n250 ) );
  NANDN U2068 ( .B(n566), .A(key[85]), .Z(\e/n249 ) );
  NANDN U2069 ( .B(n566), .A(key[84]), .Z(\e/n248 ) );
  NANDN U2070 ( .B(n566), .A(key[83]), .Z(\e/n247 ) );
  NANDN U2071 ( .B(n566), .A(key[82]), .Z(\e/n246 ) );
  NANDN U2072 ( .B(n566), .A(key[81]), .Z(\e/n245 ) );
  NANDN U2073 ( .B(n566), .A(key[80]), .Z(\e/n244 ) );
  NANDN U2074 ( .B(n566), .A(key[79]), .Z(\e/n243 ) );
  NANDN U2075 ( .B(n566), .A(key[78]), .Z(\e/n242 ) );
  NANDN U2076 ( .B(n566), .A(key[77]), .Z(\e/n241 ) );
  NANDN U2077 ( .B(n566), .A(key[76]), .Z(\e/n240 ) );
  NANDN U2078 ( .B(n566), .A(key[75]), .Z(\e/n239 ) );
  NANDN U2079 ( .B(n566), .A(key[74]), .Z(\e/n238 ) );
  NANDN U2080 ( .B(n566), .A(key[73]), .Z(\e/n237 ) );
  NANDN U2081 ( .B(n566), .A(key[72]), .Z(\e/n236 ) );
  NANDN U2082 ( .B(n566), .A(key[71]), .Z(\e/n235 ) );
  NANDN U2083 ( .B(n566), .A(key[70]), .Z(\e/n234 ) );
  NANDN U2084 ( .B(n566), .A(key[69]), .Z(\e/n233 ) );
  NANDN U2085 ( .B(n566), .A(key[68]), .Z(\e/n232 ) );
  NANDN U2086 ( .B(n566), .A(key[67]), .Z(\e/n231 ) );
  NANDN U2087 ( .B(n566), .A(key[66]), .Z(\e/n230 ) );
  NANDN U2088 ( .B(n566), .A(key[65]), .Z(\e/n229 ) );
  NANDN U2089 ( .B(n566), .A(key[64]), .Z(\e/n228 ) );
  NANDN U2090 ( .B(n566), .A(key[63]), .Z(\e/n227 ) );
  NANDN U2091 ( .B(n566), .A(key[62]), .Z(\e/n226 ) );
  NANDN U2092 ( .B(n566), .A(key[61]), .Z(\e/n225 ) );
  NANDN U2093 ( .B(n566), .A(key[60]), .Z(\e/n224 ) );
  NANDN U2094 ( .B(n566), .A(key[59]), .Z(\e/n223 ) );
  NANDN U2095 ( .B(n566), .A(key[58]), .Z(\e/n222 ) );
  NANDN U2096 ( .B(n566), .A(key[57]), .Z(\e/n221 ) );
  NANDN U2097 ( .B(n566), .A(key[56]), .Z(\e/n220 ) );
  NANDN U2098 ( .B(n566), .A(key[55]), .Z(\e/n219 ) );
  NANDN U2099 ( .B(n566), .A(key[54]), .Z(\e/n218 ) );
  NANDN U2100 ( .B(n566), .A(key[53]), .Z(\e/n217 ) );
  NANDN U2101 ( .B(n566), .A(key[52]), .Z(\e/n216 ) );
  NANDN U2102 ( .B(n566), .A(key[51]), .Z(\e/n215 ) );
  NANDN U2103 ( .B(n566), .A(key[50]), .Z(\e/n214 ) );
  NANDN U2104 ( .B(n566), .A(key[49]), .Z(\e/n213 ) );
  NANDN U2105 ( .B(n566), .A(key[48]), .Z(\e/n212 ) );
  NANDN U2106 ( .B(n566), .A(key[47]), .Z(\e/n211 ) );
  NANDN U2107 ( .B(n566), .A(key[46]), .Z(\e/n210 ) );
  NANDN U2108 ( .B(n566), .A(key[45]), .Z(\e/n209 ) );
  NANDN U2109 ( .B(n566), .A(key[44]), .Z(\e/n208 ) );
  NANDN U2110 ( .B(n566), .A(key[43]), .Z(\e/n207 ) );
  NANDN U2111 ( .B(n566), .A(key[42]), .Z(\e/n206 ) );
  NANDN U2112 ( .B(n566), .A(key[41]), .Z(\e/n205 ) );
  NANDN U2113 ( .B(n566), .A(key[40]), .Z(\e/n204 ) );
  NANDN U2114 ( .B(n566), .A(key[39]), .Z(\e/n203 ) );
  NANDN U2115 ( .B(n566), .A(key[38]), .Z(\e/n202 ) );
  NANDN U2116 ( .B(n566), .A(key[37]), .Z(\e/n201 ) );
  NANDN U2117 ( .B(n566), .A(key[36]), .Z(\e/n200 ) );
  NANDN U2118 ( .B(n566), .A(key[35]), .Z(\e/n199 ) );
  NANDN U2119 ( .B(n566), .A(key[34]), .Z(\e/n198 ) );
  NANDN U2120 ( .B(n566), .A(key[33]), .Z(\e/n197 ) );
  NANDN U2121 ( .B(n566), .A(key[32]), .Z(\e/n196 ) );
  NANDN U2122 ( .B(n566), .A(key[7]), .Z(\e/n195 ) );
  NANDN U2123 ( .B(n566), .A(key[6]), .Z(\e/n194 ) );
  NANDN U2124 ( .B(n566), .A(key[5]), .Z(\e/n193 ) );
  NANDN U2125 ( .B(n566), .A(key[4]), .Z(\e/n192 ) );
  NANDN U2126 ( .B(n566), .A(key[3]), .Z(\e/n191 ) );
  NANDN U2127 ( .B(n566), .A(key[2]), .Z(\e/n190 ) );
  NANDN U2128 ( .B(n566), .A(key[1]), .Z(\e/n189 ) );
  NANDN U2129 ( .B(n566), .A(key[0]), .Z(\e/n188 ) );
  NANDN U2130 ( .B(n1685), .A(n1688), .Z(\e/n187 ) );
  ANDN U2131 ( .A(counter[0]), .B(n1689), .Z(n1688) );
  NANDN U2132 ( .B(n1685), .A(n1690), .Z(\e/n186 ) );
  ANDN U2133 ( .A(n7), .B(n1689), .Z(n1690) );
  AND U2134 ( .A(n1691), .B(n1692), .Z(\e/n185 ) );
  NANDN U2135 ( .B(n7), .A(counter[3]), .Z(n1692) );
  NANDN U2136 ( .B(n1685), .A(n1693), .Z(n1691) );
  ANDN U2137 ( .A(n1689), .B(n7), .Z(n1693) );
  ANDN U2138 ( .A(n1694), .B(n1695), .Z(\e/n184 ) );
  NANDN U2139 ( .B(n1685), .A(n1683), .Z(n1694) );
  ANDN U2140 ( .A(n7), .B(counter[1]), .Z(n1683) );
  NAND U2141 ( .A(n1696), .B(n1697), .Z(\e/n183 ) );
  NOR U2142 ( .A(counter[2]), .B(n1698), .Z(n1697) );
  NAND U2143 ( .A(n1701), .B(n1702), .Z(\e/n182 ) );
  NOR U2144 ( .A(counter[2]), .B(n1699), .Z(n1702) );
  AND U2145 ( .A(counter[3]), .B(counter[1]), .Z(n1699) );
  IV U2146 ( .A(counter[0]), .Z(n7) );
  NOR U2147 ( .A(n1698), .B(n1695), .Z(\e/n181 ) );
  AND U2148 ( .A(counter[3]), .B(n1689), .Z(n1695) );
  ANDN U2149 ( .A(counter[0]), .B(n1703), .Z(n1698) );
  OR U2150 ( .A(n1703), .B(counter[0]), .Z(\e/n180 ) );
  AND U2151 ( .A(\e/a/SBOX[15].sbox/t[44] ), .B(\e/a/SBOX[15].sbox/y[12] ), 
        .Z(\e/a/SBOX[15].sbox/z[9] ) );
  AND U2152 ( .A(\e/a/SBOX[15].sbox/t[41] ), .B(\e/a/SBOX[15].sbox/y[10] ), 
        .Z(\e/a/SBOX[15].sbox/z[8] ) );
  AND U2153 ( .A(\e/a/SBOX[15].sbox/t[45] ), .B(\e/a/SBOX[15].sbox/y[17] ), 
        .Z(\e/a/SBOX[15].sbox/z[7] ) );
  AND U2154 ( .A(\e/a/SBOX[15].sbox/t[42] ), .B(\e/a/SBOX[15].sbox/y[11] ), 
        .Z(\e/a/SBOX[15].sbox/z[6] ) );
  AND U2155 ( .A(\e/a/SBOX[15].sbox/t[29] ), .B(\e/a/SBOX[15].sbox/y[7] ), .Z(
        \e/a/SBOX[15].sbox/z[5] ) );
  AND U2156 ( .A(\e/a/SBOX[15].sbox/t[40] ), .B(\e/a/SBOX[15].sbox/y[1] ), .Z(
        \e/a/SBOX[15].sbox/z[4] ) );
  AND U2157 ( .A(\e/a/SBOX[15].sbox/t[43] ), .B(\e/a/SBOX[15].sbox/y[16] ), 
        .Z(\e/a/SBOX[15].sbox/z[3] ) );
  ANDN U2158 ( .A(\e/a/SBOX[15].sbox/t[33] ), .B(\e/n74 ), .Z(
        \e/a/SBOX[15].sbox/z[2] ) );
  AND U2159 ( .A(\e/a/SBOX[15].sbox/t[37] ), .B(\e/a/SBOX[15].sbox/y[6] ), .Z(
        \e/a/SBOX[15].sbox/z[1] ) );
  ANDN U2160 ( .A(\e/a/SBOX[15].sbox/t[41] ), .B(n1704), .Z(
        \e/a/SBOX[15].sbox/z[17] ) );
  ANDN U2161 ( .A(\e/a/SBOX[15].sbox/t[45] ), .B(n1705), .Z(
        \e/a/SBOX[15].sbox/z[16] ) );
  ANDN U2162 ( .A(\e/a/SBOX[15].sbox/t[42] ), .B(n1706), .Z(
        \e/a/SBOX[15].sbox/z[15] ) );
  AND U2163 ( .A(\e/a/SBOX[15].sbox/t[29] ), .B(\e/a/SBOX[15].sbox/y[2] ), .Z(
        \e/a/SBOX[15].sbox/z[14] ) );
  AND U2164 ( .A(\e/a/SBOX[15].sbox/t[40] ), .B(\e/a/SBOX[15].sbox/y[5] ), .Z(
        \e/a/SBOX[15].sbox/z[13] ) );
  ANDN U2165 ( .A(\e/a/SBOX[15].sbox/t[43] ), .B(n1707), .Z(
        \e/a/SBOX[15].sbox/z[12] ) );
  AND U2166 ( .A(\e/a/SBOX[15].sbox/t[33] ), .B(\e/a/SBOX[15].sbox/y[4] ), .Z(
        \e/a/SBOX[15].sbox/z[11] ) );
  AND U2167 ( .A(\e/a/SBOX[15].sbox/t[37] ), .B(\e/a/SBOX[15].sbox/y[3] ), .Z(
        \e/a/SBOX[15].sbox/z[10] ) );
  AND U2168 ( .A(\e/a/SBOX[15].sbox/t[44] ), .B(\e/a/SBOX[15].sbox/y[15] ), 
        .Z(\e/a/SBOX[15].sbox/z[0] ) );
  AND U2169 ( .A(\e/a/SBOX[15].sbox/y[5] ), .B(\e/a/SBOX[15].sbox/y[1] ), .Z(
        \e/a/SBOX[15].sbox/t[8] ) );
  ANDN U2170 ( .A(\e/a/SBOX[15].sbox/y[16] ), .B(n1707), .Z(
        \e/a/SBOX[15].sbox/t[7] ) );
  XNOR U2171 ( .A(\e/w[3][1] ), .B(\e/w[3][7] ), .Z(n1707) );
  AND U2172 ( .A(key[97]), .B(n1687), .Z(\e/w[3][1] ) );
  ANDN U2173 ( .A(\e/a/SBOX[15].sbox/y[4] ), .B(\e/n74 ), .Z(
        \e/a/SBOX[15].sbox/t[5] ) );
  IV U2174 ( .A(\e/w[3][0] ), .Z(\e/n74 ) );
  AND U2175 ( .A(key[96]), .B(n1687), .Z(\e/w[3][0] ) );
  AND U2176 ( .A(\e/a/SBOX[15].sbox/y[3] ), .B(\e/a/SBOX[15].sbox/y[6] ), .Z(
        \e/a/SBOX[15].sbox/t[3] ) );
  AND U2177 ( .A(\e/a/SBOX[15].sbox/t[38] ), .B(\e/a/SBOX[15].sbox/t[29] ), 
        .Z(\e/a/SBOX[15].sbox/t[39] ) );
  AND U2178 ( .A(\e/a/SBOX[15].sbox/t[24] ), .B(n1708), .Z(
        \e/a/SBOX[15].sbox/t[36] ) );
  XOR U2179 ( .A(\e/a/SBOX[15].sbox/t[32] ), .B(\e/a/SBOX[15].sbox/t[26] ), 
        .Z(n1708) );
  AND U2180 ( .A(\e/a/SBOX[15].sbox/t[31] ), .B(\e/a/SBOX[15].sbox/t[30] ), 
        .Z(\e/a/SBOX[15].sbox/t[32] ) );
  AND U2181 ( .A(\e/a/SBOX[15].sbox/y[15] ), .B(\e/a/SBOX[15].sbox/y[12] ), 
        .Z(\e/a/SBOX[15].sbox/t[2] ) );
  AND U2182 ( .A(\e/a/SBOX[15].sbox/t[27] ), .B(\e/a/SBOX[15].sbox/t[25] ), 
        .Z(\e/a/SBOX[15].sbox/t[28] ) );
  AND U2183 ( .A(\e/a/SBOX[15].sbox/t[23] ), .B(\e/a/SBOX[15].sbox/t[21] ), 
        .Z(\e/a/SBOX[15].sbox/t[26] ) );
  ANDN U2184 ( .A(\e/a/SBOX[15].sbox/y[10] ), .B(n1704), .Z(
        \e/a/SBOX[15].sbox/t[15] ) );
  XNOR U2185 ( .A(\e/w[3][2] ), .B(\e/w[3][7] ), .Z(n1704) );
  ANDN U2186 ( .A(\e/a/SBOX[15].sbox/y[17] ), .B(n1705), .Z(
        \e/a/SBOX[15].sbox/t[13] ) );
  XNOR U2187 ( .A(\e/w[3][2] ), .B(\e/w[3][4] ), .Z(n1705) );
  AND U2188 ( .A(key[98]), .B(n1687), .Z(\e/w[3][2] ) );
  ANDN U2189 ( .A(\e/a/SBOX[15].sbox/y[11] ), .B(n1706), .Z(
        \e/a/SBOX[15].sbox/t[12] ) );
  XNOR U2190 ( .A(\e/w[3][4] ), .B(\e/w[3][7] ), .Z(n1706) );
  AND U2191 ( .A(key[103]), .B(n1687), .Z(\e/w[3][7] ) );
  AND U2192 ( .A(key[100]), .B(n1687), .Z(\e/w[3][4] ) );
  AND U2193 ( .A(\e/a/SBOX[15].sbox/y[2] ), .B(\e/a/SBOX[15].sbox/y[7] ), .Z(
        \e/a/SBOX[15].sbox/t[10] ) );
  AND U2194 ( .A(\e/a/SBOX[14].sbox/t[44] ), .B(\e/a/SBOX[14].sbox/y[12] ), 
        .Z(\e/a/SBOX[14].sbox/z[9] ) );
  AND U2195 ( .A(\e/a/SBOX[14].sbox/t[41] ), .B(\e/a/SBOX[14].sbox/y[10] ), 
        .Z(\e/a/SBOX[14].sbox/z[8] ) );
  AND U2196 ( .A(\e/a/SBOX[14].sbox/t[45] ), .B(\e/a/SBOX[14].sbox/y[17] ), 
        .Z(\e/a/SBOX[14].sbox/z[7] ) );
  AND U2197 ( .A(\e/a/SBOX[14].sbox/t[42] ), .B(\e/a/SBOX[14].sbox/y[11] ), 
        .Z(\e/a/SBOX[14].sbox/z[6] ) );
  AND U2198 ( .A(\e/a/SBOX[14].sbox/t[29] ), .B(\e/a/SBOX[14].sbox/y[7] ), .Z(
        \e/a/SBOX[14].sbox/z[5] ) );
  AND U2199 ( .A(\e/a/SBOX[14].sbox/t[40] ), .B(\e/a/SBOX[14].sbox/y[1] ), .Z(
        \e/a/SBOX[14].sbox/z[4] ) );
  AND U2200 ( .A(\e/a/SBOX[14].sbox/t[43] ), .B(\e/a/SBOX[14].sbox/y[16] ), 
        .Z(\e/a/SBOX[14].sbox/z[3] ) );
  ANDN U2201 ( .A(\e/a/SBOX[14].sbox/t[33] ), .B(\e/n50 ), .Z(
        \e/a/SBOX[14].sbox/z[2] ) );
  AND U2202 ( .A(\e/a/SBOX[14].sbox/t[37] ), .B(\e/a/SBOX[14].sbox/y[6] ), .Z(
        \e/a/SBOX[14].sbox/z[1] ) );
  ANDN U2203 ( .A(\e/a/SBOX[14].sbox/t[41] ), .B(n1709), .Z(
        \e/a/SBOX[14].sbox/z[17] ) );
  ANDN U2204 ( .A(\e/a/SBOX[14].sbox/t[45] ), .B(n1710), .Z(
        \e/a/SBOX[14].sbox/z[16] ) );
  ANDN U2205 ( .A(\e/a/SBOX[14].sbox/t[42] ), .B(n1711), .Z(
        \e/a/SBOX[14].sbox/z[15] ) );
  AND U2206 ( .A(\e/a/SBOX[14].sbox/t[29] ), .B(\e/a/SBOX[14].sbox/y[2] ), .Z(
        \e/a/SBOX[14].sbox/z[14] ) );
  AND U2207 ( .A(\e/a/SBOX[14].sbox/t[40] ), .B(\e/a/SBOX[14].sbox/y[5] ), .Z(
        \e/a/SBOX[14].sbox/z[13] ) );
  ANDN U2208 ( .A(\e/a/SBOX[14].sbox/t[43] ), .B(n1712), .Z(
        \e/a/SBOX[14].sbox/z[12] ) );
  AND U2209 ( .A(\e/a/SBOX[14].sbox/t[33] ), .B(\e/a/SBOX[14].sbox/y[4] ), .Z(
        \e/a/SBOX[14].sbox/z[11] ) );
  AND U2210 ( .A(\e/a/SBOX[14].sbox/t[37] ), .B(\e/a/SBOX[14].sbox/y[3] ), .Z(
        \e/a/SBOX[14].sbox/z[10] ) );
  AND U2211 ( .A(\e/a/SBOX[14].sbox/t[44] ), .B(\e/a/SBOX[14].sbox/y[15] ), 
        .Z(\e/a/SBOX[14].sbox/z[0] ) );
  AND U2212 ( .A(\e/a/SBOX[14].sbox/y[5] ), .B(\e/a/SBOX[14].sbox/y[1] ), .Z(
        \e/a/SBOX[14].sbox/t[8] ) );
  ANDN U2213 ( .A(\e/a/SBOX[14].sbox/y[16] ), .B(n1712), .Z(
        \e/a/SBOX[14].sbox/t[7] ) );
  XNOR U2214 ( .A(\e/w[3][25] ), .B(\e/w[3][31] ), .Z(n1712) );
  AND U2215 ( .A(key[121]), .B(n1687), .Z(\e/w[3][25] ) );
  ANDN U2216 ( .A(\e/a/SBOX[14].sbox/y[4] ), .B(\e/n50 ), .Z(
        \e/a/SBOX[14].sbox/t[5] ) );
  IV U2217 ( .A(\e/w[3][24] ), .Z(\e/n50 ) );
  AND U2218 ( .A(key[120]), .B(n1687), .Z(\e/w[3][24] ) );
  AND U2219 ( .A(\e/a/SBOX[14].sbox/y[3] ), .B(\e/a/SBOX[14].sbox/y[6] ), .Z(
        \e/a/SBOX[14].sbox/t[3] ) );
  AND U2220 ( .A(\e/a/SBOX[14].sbox/t[38] ), .B(\e/a/SBOX[14].sbox/t[29] ), 
        .Z(\e/a/SBOX[14].sbox/t[39] ) );
  AND U2221 ( .A(\e/a/SBOX[14].sbox/t[24] ), .B(n1713), .Z(
        \e/a/SBOX[14].sbox/t[36] ) );
  XOR U2222 ( .A(\e/a/SBOX[14].sbox/t[32] ), .B(\e/a/SBOX[14].sbox/t[26] ), 
        .Z(n1713) );
  AND U2223 ( .A(\e/a/SBOX[14].sbox/t[31] ), .B(\e/a/SBOX[14].sbox/t[30] ), 
        .Z(\e/a/SBOX[14].sbox/t[32] ) );
  AND U2224 ( .A(\e/a/SBOX[14].sbox/y[15] ), .B(\e/a/SBOX[14].sbox/y[12] ), 
        .Z(\e/a/SBOX[14].sbox/t[2] ) );
  AND U2225 ( .A(\e/a/SBOX[14].sbox/t[27] ), .B(\e/a/SBOX[14].sbox/t[25] ), 
        .Z(\e/a/SBOX[14].sbox/t[28] ) );
  AND U2226 ( .A(\e/a/SBOX[14].sbox/t[23] ), .B(\e/a/SBOX[14].sbox/t[21] ), 
        .Z(\e/a/SBOX[14].sbox/t[26] ) );
  ANDN U2227 ( .A(\e/a/SBOX[14].sbox/y[10] ), .B(n1709), .Z(
        \e/a/SBOX[14].sbox/t[15] ) );
  XNOR U2228 ( .A(\e/w[3][26] ), .B(\e/w[3][31] ), .Z(n1709) );
  ANDN U2229 ( .A(\e/a/SBOX[14].sbox/y[17] ), .B(n1710), .Z(
        \e/a/SBOX[14].sbox/t[13] ) );
  XNOR U2230 ( .A(\e/w[3][26] ), .B(\e/w[3][28] ), .Z(n1710) );
  AND U2231 ( .A(key[122]), .B(n1687), .Z(\e/w[3][26] ) );
  ANDN U2232 ( .A(\e/a/SBOX[14].sbox/y[11] ), .B(n1711), .Z(
        \e/a/SBOX[14].sbox/t[12] ) );
  XNOR U2233 ( .A(\e/w[3][28] ), .B(\e/w[3][31] ), .Z(n1711) );
  AND U2234 ( .A(key[127]), .B(n1687), .Z(\e/w[3][31] ) );
  AND U2235 ( .A(key[124]), .B(n1687), .Z(\e/w[3][28] ) );
  AND U2236 ( .A(\e/a/SBOX[14].sbox/y[2] ), .B(\e/a/SBOX[14].sbox/y[7] ), .Z(
        \e/a/SBOX[14].sbox/t[10] ) );
  AND U2237 ( .A(\e/a/SBOX[13].sbox/t[44] ), .B(\e/a/SBOX[13].sbox/y[12] ), 
        .Z(\e/a/SBOX[13].sbox/z[9] ) );
  AND U2238 ( .A(\e/a/SBOX[13].sbox/t[41] ), .B(\e/a/SBOX[13].sbox/y[10] ), 
        .Z(\e/a/SBOX[13].sbox/z[8] ) );
  AND U2239 ( .A(\e/a/SBOX[13].sbox/t[45] ), .B(\e/a/SBOX[13].sbox/y[17] ), 
        .Z(\e/a/SBOX[13].sbox/z[7] ) );
  AND U2240 ( .A(\e/a/SBOX[13].sbox/t[42] ), .B(\e/a/SBOX[13].sbox/y[11] ), 
        .Z(\e/a/SBOX[13].sbox/z[6] ) );
  AND U2241 ( .A(\e/a/SBOX[13].sbox/t[29] ), .B(\e/a/SBOX[13].sbox/y[7] ), .Z(
        \e/a/SBOX[13].sbox/z[5] ) );
  AND U2242 ( .A(\e/a/SBOX[13].sbox/t[40] ), .B(\e/a/SBOX[13].sbox/y[1] ), .Z(
        \e/a/SBOX[13].sbox/z[4] ) );
  AND U2243 ( .A(\e/a/SBOX[13].sbox/t[43] ), .B(\e/a/SBOX[13].sbox/y[16] ), 
        .Z(\e/a/SBOX[13].sbox/z[3] ) );
  ANDN U2244 ( .A(\e/a/SBOX[13].sbox/t[33] ), .B(\e/n58 ), .Z(
        \e/a/SBOX[13].sbox/z[2] ) );
  AND U2245 ( .A(\e/a/SBOX[13].sbox/t[37] ), .B(\e/a/SBOX[13].sbox/y[6] ), .Z(
        \e/a/SBOX[13].sbox/z[1] ) );
  ANDN U2246 ( .A(\e/a/SBOX[13].sbox/t[41] ), .B(n1714), .Z(
        \e/a/SBOX[13].sbox/z[17] ) );
  ANDN U2247 ( .A(\e/a/SBOX[13].sbox/t[45] ), .B(n1715), .Z(
        \e/a/SBOX[13].sbox/z[16] ) );
  ANDN U2248 ( .A(\e/a/SBOX[13].sbox/t[42] ), .B(n1716), .Z(
        \e/a/SBOX[13].sbox/z[15] ) );
  AND U2249 ( .A(\e/a/SBOX[13].sbox/t[29] ), .B(\e/a/SBOX[13].sbox/y[2] ), .Z(
        \e/a/SBOX[13].sbox/z[14] ) );
  AND U2250 ( .A(\e/a/SBOX[13].sbox/t[40] ), .B(\e/a/SBOX[13].sbox/y[5] ), .Z(
        \e/a/SBOX[13].sbox/z[13] ) );
  ANDN U2251 ( .A(\e/a/SBOX[13].sbox/t[43] ), .B(n1717), .Z(
        \e/a/SBOX[13].sbox/z[12] ) );
  AND U2252 ( .A(\e/a/SBOX[13].sbox/t[33] ), .B(\e/a/SBOX[13].sbox/y[4] ), .Z(
        \e/a/SBOX[13].sbox/z[11] ) );
  AND U2253 ( .A(\e/a/SBOX[13].sbox/t[37] ), .B(\e/a/SBOX[13].sbox/y[3] ), .Z(
        \e/a/SBOX[13].sbox/z[10] ) );
  AND U2254 ( .A(\e/a/SBOX[13].sbox/t[44] ), .B(\e/a/SBOX[13].sbox/y[15] ), 
        .Z(\e/a/SBOX[13].sbox/z[0] ) );
  AND U2255 ( .A(\e/a/SBOX[13].sbox/y[5] ), .B(\e/a/SBOX[13].sbox/y[1] ), .Z(
        \e/a/SBOX[13].sbox/t[8] ) );
  ANDN U2256 ( .A(\e/a/SBOX[13].sbox/y[16] ), .B(n1717), .Z(
        \e/a/SBOX[13].sbox/t[7] ) );
  XNOR U2257 ( .A(\e/w[3][17] ), .B(\e/w[3][23] ), .Z(n1717) );
  AND U2258 ( .A(key[113]), .B(n1687), .Z(\e/w[3][17] ) );
  ANDN U2259 ( .A(\e/a/SBOX[13].sbox/y[4] ), .B(\e/n58 ), .Z(
        \e/a/SBOX[13].sbox/t[5] ) );
  IV U2260 ( .A(\e/w[3][16] ), .Z(\e/n58 ) );
  AND U2261 ( .A(key[112]), .B(n1687), .Z(\e/w[3][16] ) );
  AND U2262 ( .A(\e/a/SBOX[13].sbox/y[3] ), .B(\e/a/SBOX[13].sbox/y[6] ), .Z(
        \e/a/SBOX[13].sbox/t[3] ) );
  AND U2263 ( .A(\e/a/SBOX[13].sbox/t[38] ), .B(\e/a/SBOX[13].sbox/t[29] ), 
        .Z(\e/a/SBOX[13].sbox/t[39] ) );
  AND U2264 ( .A(\e/a/SBOX[13].sbox/t[24] ), .B(n1718), .Z(
        \e/a/SBOX[13].sbox/t[36] ) );
  XOR U2265 ( .A(\e/a/SBOX[13].sbox/t[32] ), .B(\e/a/SBOX[13].sbox/t[26] ), 
        .Z(n1718) );
  AND U2266 ( .A(\e/a/SBOX[13].sbox/t[31] ), .B(\e/a/SBOX[13].sbox/t[30] ), 
        .Z(\e/a/SBOX[13].sbox/t[32] ) );
  AND U2267 ( .A(\e/a/SBOX[13].sbox/y[15] ), .B(\e/a/SBOX[13].sbox/y[12] ), 
        .Z(\e/a/SBOX[13].sbox/t[2] ) );
  AND U2268 ( .A(\e/a/SBOX[13].sbox/t[27] ), .B(\e/a/SBOX[13].sbox/t[25] ), 
        .Z(\e/a/SBOX[13].sbox/t[28] ) );
  AND U2269 ( .A(\e/a/SBOX[13].sbox/t[23] ), .B(\e/a/SBOX[13].sbox/t[21] ), 
        .Z(\e/a/SBOX[13].sbox/t[26] ) );
  ANDN U2270 ( .A(\e/a/SBOX[13].sbox/y[10] ), .B(n1714), .Z(
        \e/a/SBOX[13].sbox/t[15] ) );
  XNOR U2271 ( .A(\e/w[3][18] ), .B(\e/w[3][23] ), .Z(n1714) );
  ANDN U2272 ( .A(\e/a/SBOX[13].sbox/y[17] ), .B(n1715), .Z(
        \e/a/SBOX[13].sbox/t[13] ) );
  XNOR U2273 ( .A(\e/w[3][18] ), .B(\e/w[3][20] ), .Z(n1715) );
  AND U2274 ( .A(key[114]), .B(n1687), .Z(\e/w[3][18] ) );
  ANDN U2275 ( .A(\e/a/SBOX[13].sbox/y[11] ), .B(n1716), .Z(
        \e/a/SBOX[13].sbox/t[12] ) );
  XNOR U2276 ( .A(\e/w[3][20] ), .B(\e/w[3][23] ), .Z(n1716) );
  AND U2277 ( .A(key[119]), .B(n1687), .Z(\e/w[3][23] ) );
  AND U2278 ( .A(key[116]), .B(n1687), .Z(\e/w[3][20] ) );
  AND U2279 ( .A(\e/a/SBOX[13].sbox/y[2] ), .B(\e/a/SBOX[13].sbox/y[7] ), .Z(
        \e/a/SBOX[13].sbox/t[10] ) );
  AND U2280 ( .A(\e/a/SBOX[12].sbox/t[44] ), .B(\e/a/SBOX[12].sbox/y[12] ), 
        .Z(\e/a/SBOX[12].sbox/z[9] ) );
  AND U2281 ( .A(\e/a/SBOX[12].sbox/t[41] ), .B(\e/a/SBOX[12].sbox/y[10] ), 
        .Z(\e/a/SBOX[12].sbox/z[8] ) );
  AND U2282 ( .A(\e/a/SBOX[12].sbox/t[45] ), .B(\e/a/SBOX[12].sbox/y[17] ), 
        .Z(\e/a/SBOX[12].sbox/z[7] ) );
  AND U2283 ( .A(\e/a/SBOX[12].sbox/t[42] ), .B(\e/a/SBOX[12].sbox/y[11] ), 
        .Z(\e/a/SBOX[12].sbox/z[6] ) );
  AND U2284 ( .A(\e/a/SBOX[12].sbox/t[29] ), .B(\e/a/SBOX[12].sbox/y[7] ), .Z(
        \e/a/SBOX[12].sbox/z[5] ) );
  AND U2285 ( .A(\e/a/SBOX[12].sbox/t[40] ), .B(\e/a/SBOX[12].sbox/y[1] ), .Z(
        \e/a/SBOX[12].sbox/z[4] ) );
  AND U2286 ( .A(\e/a/SBOX[12].sbox/t[43] ), .B(\e/a/SBOX[12].sbox/y[16] ), 
        .Z(\e/a/SBOX[12].sbox/z[3] ) );
  ANDN U2287 ( .A(\e/a/SBOX[12].sbox/t[33] ), .B(\e/n66 ), .Z(
        \e/a/SBOX[12].sbox/z[2] ) );
  AND U2288 ( .A(\e/a/SBOX[12].sbox/t[37] ), .B(\e/a/SBOX[12].sbox/y[6] ), .Z(
        \e/a/SBOX[12].sbox/z[1] ) );
  ANDN U2289 ( .A(\e/a/SBOX[12].sbox/t[41] ), .B(n1719), .Z(
        \e/a/SBOX[12].sbox/z[17] ) );
  ANDN U2290 ( .A(\e/a/SBOX[12].sbox/t[45] ), .B(n1720), .Z(
        \e/a/SBOX[12].sbox/z[16] ) );
  ANDN U2291 ( .A(\e/a/SBOX[12].sbox/t[42] ), .B(n1721), .Z(
        \e/a/SBOX[12].sbox/z[15] ) );
  AND U2292 ( .A(\e/a/SBOX[12].sbox/t[29] ), .B(\e/a/SBOX[12].sbox/y[2] ), .Z(
        \e/a/SBOX[12].sbox/z[14] ) );
  AND U2293 ( .A(\e/a/SBOX[12].sbox/t[40] ), .B(\e/a/SBOX[12].sbox/y[5] ), .Z(
        \e/a/SBOX[12].sbox/z[13] ) );
  ANDN U2294 ( .A(\e/a/SBOX[12].sbox/t[43] ), .B(n1722), .Z(
        \e/a/SBOX[12].sbox/z[12] ) );
  AND U2295 ( .A(\e/a/SBOX[12].sbox/t[33] ), .B(\e/a/SBOX[12].sbox/y[4] ), .Z(
        \e/a/SBOX[12].sbox/z[11] ) );
  AND U2296 ( .A(\e/a/SBOX[12].sbox/t[37] ), .B(\e/a/SBOX[12].sbox/y[3] ), .Z(
        \e/a/SBOX[12].sbox/z[10] ) );
  AND U2297 ( .A(\e/a/SBOX[12].sbox/t[44] ), .B(\e/a/SBOX[12].sbox/y[15] ), 
        .Z(\e/a/SBOX[12].sbox/z[0] ) );
  AND U2298 ( .A(\e/a/SBOX[12].sbox/y[5] ), .B(\e/a/SBOX[12].sbox/y[1] ), .Z(
        \e/a/SBOX[12].sbox/t[8] ) );
  ANDN U2299 ( .A(\e/a/SBOX[12].sbox/y[16] ), .B(n1722), .Z(
        \e/a/SBOX[12].sbox/t[7] ) );
  XNOR U2300 ( .A(\e/w[3][15] ), .B(\e/w[3][9] ), .Z(n1722) );
  AND U2301 ( .A(key[105]), .B(n1687), .Z(\e/w[3][9] ) );
  ANDN U2302 ( .A(\e/a/SBOX[12].sbox/y[4] ), .B(\e/n66 ), .Z(
        \e/a/SBOX[12].sbox/t[5] ) );
  IV U2303 ( .A(\e/w[3][8] ), .Z(\e/n66 ) );
  AND U2304 ( .A(key[104]), .B(n1687), .Z(\e/w[3][8] ) );
  AND U2305 ( .A(\e/a/SBOX[12].sbox/y[3] ), .B(\e/a/SBOX[12].sbox/y[6] ), .Z(
        \e/a/SBOX[12].sbox/t[3] ) );
  AND U2306 ( .A(\e/a/SBOX[12].sbox/t[38] ), .B(\e/a/SBOX[12].sbox/t[29] ), 
        .Z(\e/a/SBOX[12].sbox/t[39] ) );
  AND U2307 ( .A(\e/a/SBOX[12].sbox/t[24] ), .B(n1723), .Z(
        \e/a/SBOX[12].sbox/t[36] ) );
  XOR U2308 ( .A(\e/a/SBOX[12].sbox/t[32] ), .B(\e/a/SBOX[12].sbox/t[26] ), 
        .Z(n1723) );
  AND U2309 ( .A(\e/a/SBOX[12].sbox/t[31] ), .B(\e/a/SBOX[12].sbox/t[30] ), 
        .Z(\e/a/SBOX[12].sbox/t[32] ) );
  AND U2310 ( .A(\e/a/SBOX[12].sbox/y[15] ), .B(\e/a/SBOX[12].sbox/y[12] ), 
        .Z(\e/a/SBOX[12].sbox/t[2] ) );
  AND U2311 ( .A(\e/a/SBOX[12].sbox/t[27] ), .B(\e/a/SBOX[12].sbox/t[25] ), 
        .Z(\e/a/SBOX[12].sbox/t[28] ) );
  AND U2312 ( .A(\e/a/SBOX[12].sbox/t[23] ), .B(\e/a/SBOX[12].sbox/t[21] ), 
        .Z(\e/a/SBOX[12].sbox/t[26] ) );
  ANDN U2313 ( .A(\e/a/SBOX[12].sbox/y[10] ), .B(n1719), .Z(
        \e/a/SBOX[12].sbox/t[15] ) );
  XNOR U2314 ( .A(\e/w[3][10] ), .B(\e/w[3][15] ), .Z(n1719) );
  ANDN U2315 ( .A(\e/a/SBOX[12].sbox/y[17] ), .B(n1720), .Z(
        \e/a/SBOX[12].sbox/t[13] ) );
  XNOR U2316 ( .A(\e/w[3][10] ), .B(\e/w[3][12] ), .Z(n1720) );
  AND U2317 ( .A(key[106]), .B(n1687), .Z(\e/w[3][10] ) );
  ANDN U2318 ( .A(\e/a/SBOX[12].sbox/y[11] ), .B(n1721), .Z(
        \e/a/SBOX[12].sbox/t[12] ) );
  XNOR U2319 ( .A(\e/w[3][12] ), .B(\e/w[3][15] ), .Z(n1721) );
  AND U2320 ( .A(key[111]), .B(n1687), .Z(\e/w[3][15] ) );
  AND U2321 ( .A(key[108]), .B(n1687), .Z(\e/w[3][12] ) );
  IV U2322 ( .A(n566), .Z(n1687) );
  AND U2323 ( .A(n1703), .B(counter[3]), .Z(n566) );
  NANDN U2324 ( .B(counter[1]), .A(n1685), .Z(n1703) );
  AND U2325 ( .A(\e/a/SBOX[12].sbox/y[2] ), .B(\e/a/SBOX[12].sbox/y[7] ), .Z(
        \e/a/SBOX[12].sbox/t[10] ) );
  AND U2326 ( .A(\b/SBOX[9].sbox/t[44] ), .B(\b/SBOX[9].sbox/y[12] ), .Z(
        \b/SBOX[9].sbox/z[9] ) );
  AND U2327 ( .A(\b/SBOX[9].sbox/t[41] ), .B(\b/SBOX[9].sbox/y[10] ), .Z(
        \b/SBOX[9].sbox/z[8] ) );
  AND U2328 ( .A(\b/SBOX[9].sbox/t[45] ), .B(\b/SBOX[9].sbox/y[17] ), .Z(
        \b/SBOX[9].sbox/z[7] ) );
  AND U2329 ( .A(\b/SBOX[9].sbox/t[42] ), .B(\b/SBOX[9].sbox/y[11] ), .Z(
        \b/SBOX[9].sbox/z[6] ) );
  AND U2330 ( .A(\b/SBOX[9].sbox/t[29] ), .B(\b/SBOX[9].sbox/y[7] ), .Z(
        \b/SBOX[9].sbox/z[5] ) );
  AND U2331 ( .A(\b/SBOX[9].sbox/t[40] ), .B(\b/SBOX[9].sbox/y[1] ), .Z(
        \b/SBOX[9].sbox/z[4] ) );
  AND U2332 ( .A(\b/SBOX[9].sbox/t[43] ), .B(\b/SBOX[9].sbox/y[16] ), .Z(
        \b/SBOX[9].sbox/z[3] ) );
  AND U2333 ( .A(msg[72]), .B(\b/SBOX[9].sbox/t[33] ), .Z(
        \b/SBOX[9].sbox/z[2] ) );
  AND U2334 ( .A(\b/SBOX[9].sbox/t[37] ), .B(\b/SBOX[9].sbox/y[6] ), .Z(
        \b/SBOX[9].sbox/z[1] ) );
  ANDN U2335 ( .A(\b/SBOX[9].sbox/t[41] ), .B(n1724), .Z(
        \b/SBOX[9].sbox/z[17] ) );
  ANDN U2336 ( .A(\b/SBOX[9].sbox/t[45] ), .B(n1725), .Z(
        \b/SBOX[9].sbox/z[16] ) );
  ANDN U2337 ( .A(\b/SBOX[9].sbox/t[42] ), .B(n1726), .Z(
        \b/SBOX[9].sbox/z[15] ) );
  AND U2338 ( .A(\b/SBOX[9].sbox/t[29] ), .B(\b/SBOX[9].sbox/y[2] ), .Z(
        \b/SBOX[9].sbox/z[14] ) );
  AND U2339 ( .A(\b/SBOX[9].sbox/t[40] ), .B(\b/SBOX[9].sbox/y[5] ), .Z(
        \b/SBOX[9].sbox/z[13] ) );
  ANDN U2340 ( .A(\b/SBOX[9].sbox/t[43] ), .B(n1727), .Z(
        \b/SBOX[9].sbox/z[12] ) );
  AND U2341 ( .A(\b/SBOX[9].sbox/t[33] ), .B(\b/SBOX[9].sbox/y[4] ), .Z(
        \b/SBOX[9].sbox/z[11] ) );
  AND U2342 ( .A(\b/SBOX[9].sbox/t[37] ), .B(\b/SBOX[9].sbox/y[3] ), .Z(
        \b/SBOX[9].sbox/z[10] ) );
  AND U2343 ( .A(\b/SBOX[9].sbox/t[44] ), .B(\b/SBOX[9].sbox/y[15] ), .Z(
        \b/SBOX[9].sbox/z[0] ) );
  AND U2344 ( .A(\b/SBOX[9].sbox/y[5] ), .B(\b/SBOX[9].sbox/y[1] ), .Z(
        \b/SBOX[9].sbox/t[8] ) );
  ANDN U2345 ( .A(\b/SBOX[9].sbox/y[16] ), .B(n1727), .Z(\b/SBOX[9].sbox/t[7] ) );
  XNOR U2346 ( .A(msg[73]), .B(msg[79]), .Z(n1727) );
  AND U2347 ( .A(\b/SBOX[9].sbox/y[4] ), .B(msg[72]), .Z(\b/SBOX[9].sbox/t[5] ) );
  AND U2348 ( .A(\b/SBOX[9].sbox/y[3] ), .B(\b/SBOX[9].sbox/y[6] ), .Z(
        \b/SBOX[9].sbox/t[3] ) );
  AND U2349 ( .A(\b/SBOX[9].sbox/t[38] ), .B(\b/SBOX[9].sbox/t[29] ), .Z(
        \b/SBOX[9].sbox/t[39] ) );
  AND U2350 ( .A(\b/SBOX[9].sbox/t[24] ), .B(n1728), .Z(\b/SBOX[9].sbox/t[36] ) );
  XOR U2351 ( .A(\b/SBOX[9].sbox/t[32] ), .B(\b/SBOX[9].sbox/t[26] ), .Z(n1728) );
  AND U2352 ( .A(\b/SBOX[9].sbox/t[31] ), .B(\b/SBOX[9].sbox/t[30] ), .Z(
        \b/SBOX[9].sbox/t[32] ) );
  AND U2353 ( .A(\b/SBOX[9].sbox/y[15] ), .B(\b/SBOX[9].sbox/y[12] ), .Z(
        \b/SBOX[9].sbox/t[2] ) );
  AND U2354 ( .A(\b/SBOX[9].sbox/t[27] ), .B(\b/SBOX[9].sbox/t[25] ), .Z(
        \b/SBOX[9].sbox/t[28] ) );
  AND U2355 ( .A(\b/SBOX[9].sbox/t[23] ), .B(\b/SBOX[9].sbox/t[21] ), .Z(
        \b/SBOX[9].sbox/t[26] ) );
  ANDN U2356 ( .A(\b/SBOX[9].sbox/y[10] ), .B(n1724), .Z(
        \b/SBOX[9].sbox/t[15] ) );
  XNOR U2357 ( .A(msg[74]), .B(msg[79]), .Z(n1724) );
  ANDN U2358 ( .A(\b/SBOX[9].sbox/y[17] ), .B(n1725), .Z(
        \b/SBOX[9].sbox/t[13] ) );
  XNOR U2359 ( .A(msg[74]), .B(msg[76]), .Z(n1725) );
  ANDN U2360 ( .A(\b/SBOX[9].sbox/y[11] ), .B(n1726), .Z(
        \b/SBOX[9].sbox/t[12] ) );
  XNOR U2361 ( .A(msg[76]), .B(msg[79]), .Z(n1726) );
  AND U2362 ( .A(\b/SBOX[9].sbox/y[2] ), .B(\b/SBOX[9].sbox/y[7] ), .Z(
        \b/SBOX[9].sbox/t[10] ) );
  AND U2363 ( .A(\b/SBOX[8].sbox/t[44] ), .B(\b/SBOX[8].sbox/y[12] ), .Z(
        \b/SBOX[8].sbox/z[9] ) );
  AND U2364 ( .A(\b/SBOX[8].sbox/t[41] ), .B(\b/SBOX[8].sbox/y[10] ), .Z(
        \b/SBOX[8].sbox/z[8] ) );
  AND U2365 ( .A(\b/SBOX[8].sbox/t[45] ), .B(\b/SBOX[8].sbox/y[17] ), .Z(
        \b/SBOX[8].sbox/z[7] ) );
  AND U2366 ( .A(\b/SBOX[8].sbox/t[42] ), .B(\b/SBOX[8].sbox/y[11] ), .Z(
        \b/SBOX[8].sbox/z[6] ) );
  AND U2367 ( .A(\b/SBOX[8].sbox/t[29] ), .B(\b/SBOX[8].sbox/y[7] ), .Z(
        \b/SBOX[8].sbox/z[5] ) );
  AND U2368 ( .A(\b/SBOX[8].sbox/t[40] ), .B(\b/SBOX[8].sbox/y[1] ), .Z(
        \b/SBOX[8].sbox/z[4] ) );
  AND U2369 ( .A(\b/SBOX[8].sbox/t[43] ), .B(\b/SBOX[8].sbox/y[16] ), .Z(
        \b/SBOX[8].sbox/z[3] ) );
  AND U2370 ( .A(msg[64]), .B(\b/SBOX[8].sbox/t[33] ), .Z(
        \b/SBOX[8].sbox/z[2] ) );
  AND U2371 ( .A(\b/SBOX[8].sbox/t[37] ), .B(\b/SBOX[8].sbox/y[6] ), .Z(
        \b/SBOX[8].sbox/z[1] ) );
  ANDN U2372 ( .A(\b/SBOX[8].sbox/t[41] ), .B(n1729), .Z(
        \b/SBOX[8].sbox/z[17] ) );
  ANDN U2373 ( .A(\b/SBOX[8].sbox/t[45] ), .B(n1730), .Z(
        \b/SBOX[8].sbox/z[16] ) );
  ANDN U2374 ( .A(\b/SBOX[8].sbox/t[42] ), .B(n1731), .Z(
        \b/SBOX[8].sbox/z[15] ) );
  AND U2375 ( .A(\b/SBOX[8].sbox/t[29] ), .B(\b/SBOX[8].sbox/y[2] ), .Z(
        \b/SBOX[8].sbox/z[14] ) );
  AND U2376 ( .A(\b/SBOX[8].sbox/t[40] ), .B(\b/SBOX[8].sbox/y[5] ), .Z(
        \b/SBOX[8].sbox/z[13] ) );
  ANDN U2377 ( .A(\b/SBOX[8].sbox/t[43] ), .B(n1732), .Z(
        \b/SBOX[8].sbox/z[12] ) );
  AND U2378 ( .A(\b/SBOX[8].sbox/t[33] ), .B(\b/SBOX[8].sbox/y[4] ), .Z(
        \b/SBOX[8].sbox/z[11] ) );
  AND U2379 ( .A(\b/SBOX[8].sbox/t[37] ), .B(\b/SBOX[8].sbox/y[3] ), .Z(
        \b/SBOX[8].sbox/z[10] ) );
  AND U2380 ( .A(\b/SBOX[8].sbox/t[44] ), .B(\b/SBOX[8].sbox/y[15] ), .Z(
        \b/SBOX[8].sbox/z[0] ) );
  AND U2381 ( .A(\b/SBOX[8].sbox/y[5] ), .B(\b/SBOX[8].sbox/y[1] ), .Z(
        \b/SBOX[8].sbox/t[8] ) );
  ANDN U2382 ( .A(\b/SBOX[8].sbox/y[16] ), .B(n1732), .Z(\b/SBOX[8].sbox/t[7] ) );
  XNOR U2383 ( .A(msg[65]), .B(msg[71]), .Z(n1732) );
  AND U2384 ( .A(\b/SBOX[8].sbox/y[4] ), .B(msg[64]), .Z(\b/SBOX[8].sbox/t[5] ) );
  AND U2385 ( .A(\b/SBOX[8].sbox/y[3] ), .B(\b/SBOX[8].sbox/y[6] ), .Z(
        \b/SBOX[8].sbox/t[3] ) );
  AND U2386 ( .A(\b/SBOX[8].sbox/t[38] ), .B(\b/SBOX[8].sbox/t[29] ), .Z(
        \b/SBOX[8].sbox/t[39] ) );
  AND U2387 ( .A(\b/SBOX[8].sbox/t[24] ), .B(n1733), .Z(\b/SBOX[8].sbox/t[36] ) );
  XOR U2388 ( .A(\b/SBOX[8].sbox/t[32] ), .B(\b/SBOX[8].sbox/t[26] ), .Z(n1733) );
  AND U2389 ( .A(\b/SBOX[8].sbox/t[31] ), .B(\b/SBOX[8].sbox/t[30] ), .Z(
        \b/SBOX[8].sbox/t[32] ) );
  AND U2390 ( .A(\b/SBOX[8].sbox/y[15] ), .B(\b/SBOX[8].sbox/y[12] ), .Z(
        \b/SBOX[8].sbox/t[2] ) );
  AND U2391 ( .A(\b/SBOX[8].sbox/t[27] ), .B(\b/SBOX[8].sbox/t[25] ), .Z(
        \b/SBOX[8].sbox/t[28] ) );
  AND U2392 ( .A(\b/SBOX[8].sbox/t[23] ), .B(\b/SBOX[8].sbox/t[21] ), .Z(
        \b/SBOX[8].sbox/t[26] ) );
  ANDN U2393 ( .A(\b/SBOX[8].sbox/y[10] ), .B(n1729), .Z(
        \b/SBOX[8].sbox/t[15] ) );
  XNOR U2394 ( .A(msg[66]), .B(msg[71]), .Z(n1729) );
  ANDN U2395 ( .A(\b/SBOX[8].sbox/y[17] ), .B(n1730), .Z(
        \b/SBOX[8].sbox/t[13] ) );
  XNOR U2396 ( .A(msg[66]), .B(msg[68]), .Z(n1730) );
  ANDN U2397 ( .A(\b/SBOX[8].sbox/y[11] ), .B(n1731), .Z(
        \b/SBOX[8].sbox/t[12] ) );
  XNOR U2398 ( .A(msg[68]), .B(msg[71]), .Z(n1731) );
  AND U2399 ( .A(\b/SBOX[8].sbox/y[2] ), .B(\b/SBOX[8].sbox/y[7] ), .Z(
        \b/SBOX[8].sbox/t[10] ) );
  AND U2400 ( .A(\b/SBOX[7].sbox/t[44] ), .B(\b/SBOX[7].sbox/y[12] ), .Z(
        \b/SBOX[7].sbox/z[9] ) );
  AND U2401 ( .A(\b/SBOX[7].sbox/t[41] ), .B(\b/SBOX[7].sbox/y[10] ), .Z(
        \b/SBOX[7].sbox/z[8] ) );
  AND U2402 ( .A(\b/SBOX[7].sbox/t[45] ), .B(\b/SBOX[7].sbox/y[17] ), .Z(
        \b/SBOX[7].sbox/z[7] ) );
  AND U2403 ( .A(\b/SBOX[7].sbox/t[42] ), .B(\b/SBOX[7].sbox/y[11] ), .Z(
        \b/SBOX[7].sbox/z[6] ) );
  AND U2404 ( .A(\b/SBOX[7].sbox/t[29] ), .B(\b/SBOX[7].sbox/y[7] ), .Z(
        \b/SBOX[7].sbox/z[5] ) );
  AND U2405 ( .A(\b/SBOX[7].sbox/t[40] ), .B(\b/SBOX[7].sbox/y[1] ), .Z(
        \b/SBOX[7].sbox/z[4] ) );
  AND U2406 ( .A(\b/SBOX[7].sbox/t[43] ), .B(\b/SBOX[7].sbox/y[16] ), .Z(
        \b/SBOX[7].sbox/z[3] ) );
  AND U2407 ( .A(msg[56]), .B(\b/SBOX[7].sbox/t[33] ), .Z(
        \b/SBOX[7].sbox/z[2] ) );
  AND U2408 ( .A(\b/SBOX[7].sbox/t[37] ), .B(\b/SBOX[7].sbox/y[6] ), .Z(
        \b/SBOX[7].sbox/z[1] ) );
  ANDN U2409 ( .A(\b/SBOX[7].sbox/t[41] ), .B(n1734), .Z(
        \b/SBOX[7].sbox/z[17] ) );
  ANDN U2410 ( .A(\b/SBOX[7].sbox/t[45] ), .B(n1735), .Z(
        \b/SBOX[7].sbox/z[16] ) );
  ANDN U2411 ( .A(\b/SBOX[7].sbox/t[42] ), .B(n1736), .Z(
        \b/SBOX[7].sbox/z[15] ) );
  AND U2412 ( .A(\b/SBOX[7].sbox/t[29] ), .B(\b/SBOX[7].sbox/y[2] ), .Z(
        \b/SBOX[7].sbox/z[14] ) );
  AND U2413 ( .A(\b/SBOX[7].sbox/t[40] ), .B(\b/SBOX[7].sbox/y[5] ), .Z(
        \b/SBOX[7].sbox/z[13] ) );
  ANDN U2414 ( .A(\b/SBOX[7].sbox/t[43] ), .B(n1737), .Z(
        \b/SBOX[7].sbox/z[12] ) );
  AND U2415 ( .A(\b/SBOX[7].sbox/t[33] ), .B(\b/SBOX[7].sbox/y[4] ), .Z(
        \b/SBOX[7].sbox/z[11] ) );
  AND U2416 ( .A(\b/SBOX[7].sbox/t[37] ), .B(\b/SBOX[7].sbox/y[3] ), .Z(
        \b/SBOX[7].sbox/z[10] ) );
  AND U2417 ( .A(\b/SBOX[7].sbox/t[44] ), .B(\b/SBOX[7].sbox/y[15] ), .Z(
        \b/SBOX[7].sbox/z[0] ) );
  AND U2418 ( .A(\b/SBOX[7].sbox/y[5] ), .B(\b/SBOX[7].sbox/y[1] ), .Z(
        \b/SBOX[7].sbox/t[8] ) );
  ANDN U2419 ( .A(\b/SBOX[7].sbox/y[16] ), .B(n1737), .Z(\b/SBOX[7].sbox/t[7] ) );
  XNOR U2420 ( .A(msg[57]), .B(msg[63]), .Z(n1737) );
  AND U2421 ( .A(\b/SBOX[7].sbox/y[4] ), .B(msg[56]), .Z(\b/SBOX[7].sbox/t[5] ) );
  AND U2422 ( .A(\b/SBOX[7].sbox/y[3] ), .B(\b/SBOX[7].sbox/y[6] ), .Z(
        \b/SBOX[7].sbox/t[3] ) );
  AND U2423 ( .A(\b/SBOX[7].sbox/t[38] ), .B(\b/SBOX[7].sbox/t[29] ), .Z(
        \b/SBOX[7].sbox/t[39] ) );
  AND U2424 ( .A(\b/SBOX[7].sbox/t[24] ), .B(n1738), .Z(\b/SBOX[7].sbox/t[36] ) );
  XOR U2425 ( .A(\b/SBOX[7].sbox/t[32] ), .B(\b/SBOX[7].sbox/t[26] ), .Z(n1738) );
  AND U2426 ( .A(\b/SBOX[7].sbox/t[31] ), .B(\b/SBOX[7].sbox/t[30] ), .Z(
        \b/SBOX[7].sbox/t[32] ) );
  AND U2427 ( .A(\b/SBOX[7].sbox/y[15] ), .B(\b/SBOX[7].sbox/y[12] ), .Z(
        \b/SBOX[7].sbox/t[2] ) );
  AND U2428 ( .A(\b/SBOX[7].sbox/t[27] ), .B(\b/SBOX[7].sbox/t[25] ), .Z(
        \b/SBOX[7].sbox/t[28] ) );
  AND U2429 ( .A(\b/SBOX[7].sbox/t[23] ), .B(\b/SBOX[7].sbox/t[21] ), .Z(
        \b/SBOX[7].sbox/t[26] ) );
  ANDN U2430 ( .A(\b/SBOX[7].sbox/y[10] ), .B(n1734), .Z(
        \b/SBOX[7].sbox/t[15] ) );
  XNOR U2431 ( .A(msg[58]), .B(msg[63]), .Z(n1734) );
  ANDN U2432 ( .A(\b/SBOX[7].sbox/y[17] ), .B(n1735), .Z(
        \b/SBOX[7].sbox/t[13] ) );
  XNOR U2433 ( .A(msg[58]), .B(msg[60]), .Z(n1735) );
  ANDN U2434 ( .A(\b/SBOX[7].sbox/y[11] ), .B(n1736), .Z(
        \b/SBOX[7].sbox/t[12] ) );
  XNOR U2435 ( .A(msg[60]), .B(msg[63]), .Z(n1736) );
  AND U2436 ( .A(\b/SBOX[7].sbox/y[2] ), .B(\b/SBOX[7].sbox/y[7] ), .Z(
        \b/SBOX[7].sbox/t[10] ) );
  AND U2437 ( .A(\b/SBOX[6].sbox/t[44] ), .B(\b/SBOX[6].sbox/y[12] ), .Z(
        \b/SBOX[6].sbox/z[9] ) );
  AND U2438 ( .A(\b/SBOX[6].sbox/t[41] ), .B(\b/SBOX[6].sbox/y[10] ), .Z(
        \b/SBOX[6].sbox/z[8] ) );
  AND U2439 ( .A(\b/SBOX[6].sbox/t[45] ), .B(\b/SBOX[6].sbox/y[17] ), .Z(
        \b/SBOX[6].sbox/z[7] ) );
  AND U2440 ( .A(\b/SBOX[6].sbox/t[42] ), .B(\b/SBOX[6].sbox/y[11] ), .Z(
        \b/SBOX[6].sbox/z[6] ) );
  AND U2441 ( .A(\b/SBOX[6].sbox/t[29] ), .B(\b/SBOX[6].sbox/y[7] ), .Z(
        \b/SBOX[6].sbox/z[5] ) );
  AND U2442 ( .A(\b/SBOX[6].sbox/t[40] ), .B(\b/SBOX[6].sbox/y[1] ), .Z(
        \b/SBOX[6].sbox/z[4] ) );
  AND U2443 ( .A(\b/SBOX[6].sbox/t[43] ), .B(\b/SBOX[6].sbox/y[16] ), .Z(
        \b/SBOX[6].sbox/z[3] ) );
  AND U2444 ( .A(msg[48]), .B(\b/SBOX[6].sbox/t[33] ), .Z(
        \b/SBOX[6].sbox/z[2] ) );
  AND U2445 ( .A(\b/SBOX[6].sbox/t[37] ), .B(\b/SBOX[6].sbox/y[6] ), .Z(
        \b/SBOX[6].sbox/z[1] ) );
  ANDN U2446 ( .A(\b/SBOX[6].sbox/t[41] ), .B(n1739), .Z(
        \b/SBOX[6].sbox/z[17] ) );
  ANDN U2447 ( .A(\b/SBOX[6].sbox/t[45] ), .B(n1740), .Z(
        \b/SBOX[6].sbox/z[16] ) );
  ANDN U2448 ( .A(\b/SBOX[6].sbox/t[42] ), .B(n1741), .Z(
        \b/SBOX[6].sbox/z[15] ) );
  AND U2449 ( .A(\b/SBOX[6].sbox/t[29] ), .B(\b/SBOX[6].sbox/y[2] ), .Z(
        \b/SBOX[6].sbox/z[14] ) );
  AND U2450 ( .A(\b/SBOX[6].sbox/t[40] ), .B(\b/SBOX[6].sbox/y[5] ), .Z(
        \b/SBOX[6].sbox/z[13] ) );
  ANDN U2451 ( .A(\b/SBOX[6].sbox/t[43] ), .B(n1742), .Z(
        \b/SBOX[6].sbox/z[12] ) );
  AND U2452 ( .A(\b/SBOX[6].sbox/t[33] ), .B(\b/SBOX[6].sbox/y[4] ), .Z(
        \b/SBOX[6].sbox/z[11] ) );
  AND U2453 ( .A(\b/SBOX[6].sbox/t[37] ), .B(\b/SBOX[6].sbox/y[3] ), .Z(
        \b/SBOX[6].sbox/z[10] ) );
  AND U2454 ( .A(\b/SBOX[6].sbox/t[44] ), .B(\b/SBOX[6].sbox/y[15] ), .Z(
        \b/SBOX[6].sbox/z[0] ) );
  AND U2455 ( .A(\b/SBOX[6].sbox/y[5] ), .B(\b/SBOX[6].sbox/y[1] ), .Z(
        \b/SBOX[6].sbox/t[8] ) );
  ANDN U2456 ( .A(\b/SBOX[6].sbox/y[16] ), .B(n1742), .Z(\b/SBOX[6].sbox/t[7] ) );
  XNOR U2457 ( .A(msg[49]), .B(msg[55]), .Z(n1742) );
  AND U2458 ( .A(\b/SBOX[6].sbox/y[4] ), .B(msg[48]), .Z(\b/SBOX[6].sbox/t[5] ) );
  AND U2459 ( .A(\b/SBOX[6].sbox/y[3] ), .B(\b/SBOX[6].sbox/y[6] ), .Z(
        \b/SBOX[6].sbox/t[3] ) );
  AND U2460 ( .A(\b/SBOX[6].sbox/t[38] ), .B(\b/SBOX[6].sbox/t[29] ), .Z(
        \b/SBOX[6].sbox/t[39] ) );
  AND U2461 ( .A(\b/SBOX[6].sbox/t[24] ), .B(n1743), .Z(\b/SBOX[6].sbox/t[36] ) );
  XOR U2462 ( .A(\b/SBOX[6].sbox/t[32] ), .B(\b/SBOX[6].sbox/t[26] ), .Z(n1743) );
  AND U2463 ( .A(\b/SBOX[6].sbox/t[31] ), .B(\b/SBOX[6].sbox/t[30] ), .Z(
        \b/SBOX[6].sbox/t[32] ) );
  AND U2464 ( .A(\b/SBOX[6].sbox/y[15] ), .B(\b/SBOX[6].sbox/y[12] ), .Z(
        \b/SBOX[6].sbox/t[2] ) );
  AND U2465 ( .A(\b/SBOX[6].sbox/t[27] ), .B(\b/SBOX[6].sbox/t[25] ), .Z(
        \b/SBOX[6].sbox/t[28] ) );
  AND U2466 ( .A(\b/SBOX[6].sbox/t[23] ), .B(\b/SBOX[6].sbox/t[21] ), .Z(
        \b/SBOX[6].sbox/t[26] ) );
  ANDN U2467 ( .A(\b/SBOX[6].sbox/y[10] ), .B(n1739), .Z(
        \b/SBOX[6].sbox/t[15] ) );
  XNOR U2468 ( .A(msg[50]), .B(msg[55]), .Z(n1739) );
  ANDN U2469 ( .A(\b/SBOX[6].sbox/y[17] ), .B(n1740), .Z(
        \b/SBOX[6].sbox/t[13] ) );
  XNOR U2470 ( .A(msg[50]), .B(msg[52]), .Z(n1740) );
  ANDN U2471 ( .A(\b/SBOX[6].sbox/y[11] ), .B(n1741), .Z(
        \b/SBOX[6].sbox/t[12] ) );
  XNOR U2472 ( .A(msg[52]), .B(msg[55]), .Z(n1741) );
  AND U2473 ( .A(\b/SBOX[6].sbox/y[2] ), .B(\b/SBOX[6].sbox/y[7] ), .Z(
        \b/SBOX[6].sbox/t[10] ) );
  AND U2474 ( .A(\b/SBOX[5].sbox/t[44] ), .B(\b/SBOX[5].sbox/y[12] ), .Z(
        \b/SBOX[5].sbox/z[9] ) );
  AND U2475 ( .A(\b/SBOX[5].sbox/t[41] ), .B(\b/SBOX[5].sbox/y[10] ), .Z(
        \b/SBOX[5].sbox/z[8] ) );
  AND U2476 ( .A(\b/SBOX[5].sbox/t[45] ), .B(\b/SBOX[5].sbox/y[17] ), .Z(
        \b/SBOX[5].sbox/z[7] ) );
  AND U2477 ( .A(\b/SBOX[5].sbox/t[42] ), .B(\b/SBOX[5].sbox/y[11] ), .Z(
        \b/SBOX[5].sbox/z[6] ) );
  AND U2478 ( .A(\b/SBOX[5].sbox/t[29] ), .B(\b/SBOX[5].sbox/y[7] ), .Z(
        \b/SBOX[5].sbox/z[5] ) );
  AND U2479 ( .A(\b/SBOX[5].sbox/t[40] ), .B(\b/SBOX[5].sbox/y[1] ), .Z(
        \b/SBOX[5].sbox/z[4] ) );
  AND U2480 ( .A(\b/SBOX[5].sbox/t[43] ), .B(\b/SBOX[5].sbox/y[16] ), .Z(
        \b/SBOX[5].sbox/z[3] ) );
  AND U2481 ( .A(msg[40]), .B(\b/SBOX[5].sbox/t[33] ), .Z(
        \b/SBOX[5].sbox/z[2] ) );
  AND U2482 ( .A(\b/SBOX[5].sbox/t[37] ), .B(\b/SBOX[5].sbox/y[6] ), .Z(
        \b/SBOX[5].sbox/z[1] ) );
  ANDN U2483 ( .A(\b/SBOX[5].sbox/t[41] ), .B(n1744), .Z(
        \b/SBOX[5].sbox/z[17] ) );
  ANDN U2484 ( .A(\b/SBOX[5].sbox/t[45] ), .B(n1745), .Z(
        \b/SBOX[5].sbox/z[16] ) );
  ANDN U2485 ( .A(\b/SBOX[5].sbox/t[42] ), .B(n1746), .Z(
        \b/SBOX[5].sbox/z[15] ) );
  AND U2486 ( .A(\b/SBOX[5].sbox/t[29] ), .B(\b/SBOX[5].sbox/y[2] ), .Z(
        \b/SBOX[5].sbox/z[14] ) );
  AND U2487 ( .A(\b/SBOX[5].sbox/t[40] ), .B(\b/SBOX[5].sbox/y[5] ), .Z(
        \b/SBOX[5].sbox/z[13] ) );
  ANDN U2488 ( .A(\b/SBOX[5].sbox/t[43] ), .B(n1747), .Z(
        \b/SBOX[5].sbox/z[12] ) );
  AND U2489 ( .A(\b/SBOX[5].sbox/t[33] ), .B(\b/SBOX[5].sbox/y[4] ), .Z(
        \b/SBOX[5].sbox/z[11] ) );
  AND U2490 ( .A(\b/SBOX[5].sbox/t[37] ), .B(\b/SBOX[5].sbox/y[3] ), .Z(
        \b/SBOX[5].sbox/z[10] ) );
  AND U2491 ( .A(\b/SBOX[5].sbox/t[44] ), .B(\b/SBOX[5].sbox/y[15] ), .Z(
        \b/SBOX[5].sbox/z[0] ) );
  AND U2492 ( .A(\b/SBOX[5].sbox/y[5] ), .B(\b/SBOX[5].sbox/y[1] ), .Z(
        \b/SBOX[5].sbox/t[8] ) );
  ANDN U2493 ( .A(\b/SBOX[5].sbox/y[16] ), .B(n1747), .Z(\b/SBOX[5].sbox/t[7] ) );
  XNOR U2494 ( .A(msg[41]), .B(msg[47]), .Z(n1747) );
  AND U2495 ( .A(\b/SBOX[5].sbox/y[4] ), .B(msg[40]), .Z(\b/SBOX[5].sbox/t[5] ) );
  AND U2496 ( .A(\b/SBOX[5].sbox/y[3] ), .B(\b/SBOX[5].sbox/y[6] ), .Z(
        \b/SBOX[5].sbox/t[3] ) );
  AND U2497 ( .A(\b/SBOX[5].sbox/t[38] ), .B(\b/SBOX[5].sbox/t[29] ), .Z(
        \b/SBOX[5].sbox/t[39] ) );
  AND U2498 ( .A(\b/SBOX[5].sbox/t[24] ), .B(n1748), .Z(\b/SBOX[5].sbox/t[36] ) );
  XOR U2499 ( .A(\b/SBOX[5].sbox/t[32] ), .B(\b/SBOX[5].sbox/t[26] ), .Z(n1748) );
  AND U2500 ( .A(\b/SBOX[5].sbox/t[31] ), .B(\b/SBOX[5].sbox/t[30] ), .Z(
        \b/SBOX[5].sbox/t[32] ) );
  AND U2501 ( .A(\b/SBOX[5].sbox/y[15] ), .B(\b/SBOX[5].sbox/y[12] ), .Z(
        \b/SBOX[5].sbox/t[2] ) );
  AND U2502 ( .A(\b/SBOX[5].sbox/t[27] ), .B(\b/SBOX[5].sbox/t[25] ), .Z(
        \b/SBOX[5].sbox/t[28] ) );
  AND U2503 ( .A(\b/SBOX[5].sbox/t[23] ), .B(\b/SBOX[5].sbox/t[21] ), .Z(
        \b/SBOX[5].sbox/t[26] ) );
  ANDN U2504 ( .A(\b/SBOX[5].sbox/y[10] ), .B(n1744), .Z(
        \b/SBOX[5].sbox/t[15] ) );
  XNOR U2505 ( .A(msg[42]), .B(msg[47]), .Z(n1744) );
  ANDN U2506 ( .A(\b/SBOX[5].sbox/y[17] ), .B(n1745), .Z(
        \b/SBOX[5].sbox/t[13] ) );
  XNOR U2507 ( .A(msg[42]), .B(msg[44]), .Z(n1745) );
  ANDN U2508 ( .A(\b/SBOX[5].sbox/y[11] ), .B(n1746), .Z(
        \b/SBOX[5].sbox/t[12] ) );
  XNOR U2509 ( .A(msg[44]), .B(msg[47]), .Z(n1746) );
  AND U2510 ( .A(\b/SBOX[5].sbox/y[2] ), .B(\b/SBOX[5].sbox/y[7] ), .Z(
        \b/SBOX[5].sbox/t[10] ) );
  AND U2511 ( .A(\b/SBOX[4].sbox/t[44] ), .B(\b/SBOX[4].sbox/y[12] ), .Z(
        \b/SBOX[4].sbox/z[9] ) );
  AND U2512 ( .A(\b/SBOX[4].sbox/t[41] ), .B(\b/SBOX[4].sbox/y[10] ), .Z(
        \b/SBOX[4].sbox/z[8] ) );
  AND U2513 ( .A(\b/SBOX[4].sbox/t[45] ), .B(\b/SBOX[4].sbox/y[17] ), .Z(
        \b/SBOX[4].sbox/z[7] ) );
  AND U2514 ( .A(\b/SBOX[4].sbox/t[42] ), .B(\b/SBOX[4].sbox/y[11] ), .Z(
        \b/SBOX[4].sbox/z[6] ) );
  AND U2515 ( .A(\b/SBOX[4].sbox/t[29] ), .B(\b/SBOX[4].sbox/y[7] ), .Z(
        \b/SBOX[4].sbox/z[5] ) );
  AND U2516 ( .A(\b/SBOX[4].sbox/t[40] ), .B(\b/SBOX[4].sbox/y[1] ), .Z(
        \b/SBOX[4].sbox/z[4] ) );
  AND U2517 ( .A(\b/SBOX[4].sbox/t[43] ), .B(\b/SBOX[4].sbox/y[16] ), .Z(
        \b/SBOX[4].sbox/z[3] ) );
  AND U2518 ( .A(msg[32]), .B(\b/SBOX[4].sbox/t[33] ), .Z(
        \b/SBOX[4].sbox/z[2] ) );
  AND U2519 ( .A(\b/SBOX[4].sbox/t[37] ), .B(\b/SBOX[4].sbox/y[6] ), .Z(
        \b/SBOX[4].sbox/z[1] ) );
  ANDN U2520 ( .A(\b/SBOX[4].sbox/t[41] ), .B(n1749), .Z(
        \b/SBOX[4].sbox/z[17] ) );
  ANDN U2521 ( .A(\b/SBOX[4].sbox/t[45] ), .B(n1750), .Z(
        \b/SBOX[4].sbox/z[16] ) );
  ANDN U2522 ( .A(\b/SBOX[4].sbox/t[42] ), .B(n1751), .Z(
        \b/SBOX[4].sbox/z[15] ) );
  AND U2523 ( .A(\b/SBOX[4].sbox/t[29] ), .B(\b/SBOX[4].sbox/y[2] ), .Z(
        \b/SBOX[4].sbox/z[14] ) );
  AND U2524 ( .A(\b/SBOX[4].sbox/t[40] ), .B(\b/SBOX[4].sbox/y[5] ), .Z(
        \b/SBOX[4].sbox/z[13] ) );
  ANDN U2525 ( .A(\b/SBOX[4].sbox/t[43] ), .B(n1752), .Z(
        \b/SBOX[4].sbox/z[12] ) );
  AND U2526 ( .A(\b/SBOX[4].sbox/t[33] ), .B(\b/SBOX[4].sbox/y[4] ), .Z(
        \b/SBOX[4].sbox/z[11] ) );
  AND U2527 ( .A(\b/SBOX[4].sbox/t[37] ), .B(\b/SBOX[4].sbox/y[3] ), .Z(
        \b/SBOX[4].sbox/z[10] ) );
  AND U2528 ( .A(\b/SBOX[4].sbox/t[44] ), .B(\b/SBOX[4].sbox/y[15] ), .Z(
        \b/SBOX[4].sbox/z[0] ) );
  AND U2529 ( .A(\b/SBOX[4].sbox/y[5] ), .B(\b/SBOX[4].sbox/y[1] ), .Z(
        \b/SBOX[4].sbox/t[8] ) );
  ANDN U2530 ( .A(\b/SBOX[4].sbox/y[16] ), .B(n1752), .Z(\b/SBOX[4].sbox/t[7] ) );
  XNOR U2531 ( .A(msg[33]), .B(msg[39]), .Z(n1752) );
  AND U2532 ( .A(\b/SBOX[4].sbox/y[4] ), .B(msg[32]), .Z(\b/SBOX[4].sbox/t[5] ) );
  AND U2533 ( .A(\b/SBOX[4].sbox/y[3] ), .B(\b/SBOX[4].sbox/y[6] ), .Z(
        \b/SBOX[4].sbox/t[3] ) );
  AND U2534 ( .A(\b/SBOX[4].sbox/t[38] ), .B(\b/SBOX[4].sbox/t[29] ), .Z(
        \b/SBOX[4].sbox/t[39] ) );
  AND U2535 ( .A(\b/SBOX[4].sbox/t[24] ), .B(n1753), .Z(\b/SBOX[4].sbox/t[36] ) );
  XOR U2536 ( .A(\b/SBOX[4].sbox/t[32] ), .B(\b/SBOX[4].sbox/t[26] ), .Z(n1753) );
  AND U2537 ( .A(\b/SBOX[4].sbox/t[31] ), .B(\b/SBOX[4].sbox/t[30] ), .Z(
        \b/SBOX[4].sbox/t[32] ) );
  AND U2538 ( .A(\b/SBOX[4].sbox/y[15] ), .B(\b/SBOX[4].sbox/y[12] ), .Z(
        \b/SBOX[4].sbox/t[2] ) );
  AND U2539 ( .A(\b/SBOX[4].sbox/t[27] ), .B(\b/SBOX[4].sbox/t[25] ), .Z(
        \b/SBOX[4].sbox/t[28] ) );
  AND U2540 ( .A(\b/SBOX[4].sbox/t[23] ), .B(\b/SBOX[4].sbox/t[21] ), .Z(
        \b/SBOX[4].sbox/t[26] ) );
  ANDN U2541 ( .A(\b/SBOX[4].sbox/y[10] ), .B(n1749), .Z(
        \b/SBOX[4].sbox/t[15] ) );
  XNOR U2542 ( .A(msg[34]), .B(msg[39]), .Z(n1749) );
  ANDN U2543 ( .A(\b/SBOX[4].sbox/y[17] ), .B(n1750), .Z(
        \b/SBOX[4].sbox/t[13] ) );
  XNOR U2544 ( .A(msg[34]), .B(msg[36]), .Z(n1750) );
  ANDN U2545 ( .A(\b/SBOX[4].sbox/y[11] ), .B(n1751), .Z(
        \b/SBOX[4].sbox/t[12] ) );
  XNOR U2546 ( .A(msg[36]), .B(msg[39]), .Z(n1751) );
  AND U2547 ( .A(\b/SBOX[4].sbox/y[2] ), .B(\b/SBOX[4].sbox/y[7] ), .Z(
        \b/SBOX[4].sbox/t[10] ) );
  AND U2548 ( .A(\b/SBOX[3].sbox/t[44] ), .B(\b/SBOX[3].sbox/y[12] ), .Z(
        \b/SBOX[3].sbox/z[9] ) );
  AND U2549 ( .A(\b/SBOX[3].sbox/t[41] ), .B(\b/SBOX[3].sbox/y[10] ), .Z(
        \b/SBOX[3].sbox/z[8] ) );
  AND U2550 ( .A(\b/SBOX[3].sbox/t[45] ), .B(\b/SBOX[3].sbox/y[17] ), .Z(
        \b/SBOX[3].sbox/z[7] ) );
  AND U2551 ( .A(\b/SBOX[3].sbox/t[42] ), .B(\b/SBOX[3].sbox/y[11] ), .Z(
        \b/SBOX[3].sbox/z[6] ) );
  AND U2552 ( .A(\b/SBOX[3].sbox/t[29] ), .B(\b/SBOX[3].sbox/y[7] ), .Z(
        \b/SBOX[3].sbox/z[5] ) );
  AND U2553 ( .A(\b/SBOX[3].sbox/t[40] ), .B(\b/SBOX[3].sbox/y[1] ), .Z(
        \b/SBOX[3].sbox/z[4] ) );
  AND U2554 ( .A(\b/SBOX[3].sbox/t[43] ), .B(\b/SBOX[3].sbox/y[16] ), .Z(
        \b/SBOX[3].sbox/z[3] ) );
  AND U2555 ( .A(msg[24]), .B(\b/SBOX[3].sbox/t[33] ), .Z(
        \b/SBOX[3].sbox/z[2] ) );
  AND U2556 ( .A(\b/SBOX[3].sbox/t[37] ), .B(\b/SBOX[3].sbox/y[6] ), .Z(
        \b/SBOX[3].sbox/z[1] ) );
  ANDN U2557 ( .A(\b/SBOX[3].sbox/t[41] ), .B(n1754), .Z(
        \b/SBOX[3].sbox/z[17] ) );
  ANDN U2558 ( .A(\b/SBOX[3].sbox/t[45] ), .B(n1755), .Z(
        \b/SBOX[3].sbox/z[16] ) );
  ANDN U2559 ( .A(\b/SBOX[3].sbox/t[42] ), .B(n1756), .Z(
        \b/SBOX[3].sbox/z[15] ) );
  AND U2560 ( .A(\b/SBOX[3].sbox/t[29] ), .B(\b/SBOX[3].sbox/y[2] ), .Z(
        \b/SBOX[3].sbox/z[14] ) );
  AND U2561 ( .A(\b/SBOX[3].sbox/t[40] ), .B(\b/SBOX[3].sbox/y[5] ), .Z(
        \b/SBOX[3].sbox/z[13] ) );
  ANDN U2562 ( .A(\b/SBOX[3].sbox/t[43] ), .B(n1757), .Z(
        \b/SBOX[3].sbox/z[12] ) );
  AND U2563 ( .A(\b/SBOX[3].sbox/t[33] ), .B(\b/SBOX[3].sbox/y[4] ), .Z(
        \b/SBOX[3].sbox/z[11] ) );
  AND U2564 ( .A(\b/SBOX[3].sbox/t[37] ), .B(\b/SBOX[3].sbox/y[3] ), .Z(
        \b/SBOX[3].sbox/z[10] ) );
  AND U2565 ( .A(\b/SBOX[3].sbox/t[44] ), .B(\b/SBOX[3].sbox/y[15] ), .Z(
        \b/SBOX[3].sbox/z[0] ) );
  AND U2566 ( .A(\b/SBOX[3].sbox/y[5] ), .B(\b/SBOX[3].sbox/y[1] ), .Z(
        \b/SBOX[3].sbox/t[8] ) );
  ANDN U2567 ( .A(\b/SBOX[3].sbox/y[16] ), .B(n1757), .Z(\b/SBOX[3].sbox/t[7] ) );
  XNOR U2568 ( .A(msg[25]), .B(msg[31]), .Z(n1757) );
  AND U2569 ( .A(\b/SBOX[3].sbox/y[4] ), .B(msg[24]), .Z(\b/SBOX[3].sbox/t[5] ) );
  AND U2570 ( .A(\b/SBOX[3].sbox/y[3] ), .B(\b/SBOX[3].sbox/y[6] ), .Z(
        \b/SBOX[3].sbox/t[3] ) );
  AND U2571 ( .A(\b/SBOX[3].sbox/t[38] ), .B(\b/SBOX[3].sbox/t[29] ), .Z(
        \b/SBOX[3].sbox/t[39] ) );
  AND U2572 ( .A(\b/SBOX[3].sbox/t[24] ), .B(n1758), .Z(\b/SBOX[3].sbox/t[36] ) );
  XOR U2573 ( .A(\b/SBOX[3].sbox/t[32] ), .B(\b/SBOX[3].sbox/t[26] ), .Z(n1758) );
  AND U2574 ( .A(\b/SBOX[3].sbox/t[31] ), .B(\b/SBOX[3].sbox/t[30] ), .Z(
        \b/SBOX[3].sbox/t[32] ) );
  AND U2575 ( .A(\b/SBOX[3].sbox/y[15] ), .B(\b/SBOX[3].sbox/y[12] ), .Z(
        \b/SBOX[3].sbox/t[2] ) );
  AND U2576 ( .A(\b/SBOX[3].sbox/t[27] ), .B(\b/SBOX[3].sbox/t[25] ), .Z(
        \b/SBOX[3].sbox/t[28] ) );
  AND U2577 ( .A(\b/SBOX[3].sbox/t[23] ), .B(\b/SBOX[3].sbox/t[21] ), .Z(
        \b/SBOX[3].sbox/t[26] ) );
  ANDN U2578 ( .A(\b/SBOX[3].sbox/y[10] ), .B(n1754), .Z(
        \b/SBOX[3].sbox/t[15] ) );
  XNOR U2579 ( .A(msg[26]), .B(msg[31]), .Z(n1754) );
  ANDN U2580 ( .A(\b/SBOX[3].sbox/y[17] ), .B(n1755), .Z(
        \b/SBOX[3].sbox/t[13] ) );
  XNOR U2581 ( .A(msg[26]), .B(msg[28]), .Z(n1755) );
  ANDN U2582 ( .A(\b/SBOX[3].sbox/y[11] ), .B(n1756), .Z(
        \b/SBOX[3].sbox/t[12] ) );
  XNOR U2583 ( .A(msg[28]), .B(msg[31]), .Z(n1756) );
  AND U2584 ( .A(\b/SBOX[3].sbox/y[2] ), .B(\b/SBOX[3].sbox/y[7] ), .Z(
        \b/SBOX[3].sbox/t[10] ) );
  AND U2585 ( .A(\b/SBOX[2].sbox/t[44] ), .B(\b/SBOX[2].sbox/y[12] ), .Z(
        \b/SBOX[2].sbox/z[9] ) );
  AND U2586 ( .A(\b/SBOX[2].sbox/t[41] ), .B(\b/SBOX[2].sbox/y[10] ), .Z(
        \b/SBOX[2].sbox/z[8] ) );
  AND U2587 ( .A(\b/SBOX[2].sbox/t[45] ), .B(\b/SBOX[2].sbox/y[17] ), .Z(
        \b/SBOX[2].sbox/z[7] ) );
  AND U2588 ( .A(\b/SBOX[2].sbox/t[42] ), .B(\b/SBOX[2].sbox/y[11] ), .Z(
        \b/SBOX[2].sbox/z[6] ) );
  AND U2589 ( .A(\b/SBOX[2].sbox/t[29] ), .B(\b/SBOX[2].sbox/y[7] ), .Z(
        \b/SBOX[2].sbox/z[5] ) );
  AND U2590 ( .A(\b/SBOX[2].sbox/t[40] ), .B(\b/SBOX[2].sbox/y[1] ), .Z(
        \b/SBOX[2].sbox/z[4] ) );
  AND U2591 ( .A(\b/SBOX[2].sbox/t[43] ), .B(\b/SBOX[2].sbox/y[16] ), .Z(
        \b/SBOX[2].sbox/z[3] ) );
  AND U2592 ( .A(msg[16]), .B(\b/SBOX[2].sbox/t[33] ), .Z(
        \b/SBOX[2].sbox/z[2] ) );
  AND U2593 ( .A(\b/SBOX[2].sbox/t[37] ), .B(\b/SBOX[2].sbox/y[6] ), .Z(
        \b/SBOX[2].sbox/z[1] ) );
  ANDN U2594 ( .A(\b/SBOX[2].sbox/t[41] ), .B(n1759), .Z(
        \b/SBOX[2].sbox/z[17] ) );
  ANDN U2595 ( .A(\b/SBOX[2].sbox/t[45] ), .B(n1760), .Z(
        \b/SBOX[2].sbox/z[16] ) );
  ANDN U2596 ( .A(\b/SBOX[2].sbox/t[42] ), .B(n1761), .Z(
        \b/SBOX[2].sbox/z[15] ) );
  AND U2597 ( .A(\b/SBOX[2].sbox/t[29] ), .B(\b/SBOX[2].sbox/y[2] ), .Z(
        \b/SBOX[2].sbox/z[14] ) );
  AND U2598 ( .A(\b/SBOX[2].sbox/t[40] ), .B(\b/SBOX[2].sbox/y[5] ), .Z(
        \b/SBOX[2].sbox/z[13] ) );
  ANDN U2599 ( .A(\b/SBOX[2].sbox/t[43] ), .B(n1762), .Z(
        \b/SBOX[2].sbox/z[12] ) );
  AND U2600 ( .A(\b/SBOX[2].sbox/t[33] ), .B(\b/SBOX[2].sbox/y[4] ), .Z(
        \b/SBOX[2].sbox/z[11] ) );
  AND U2601 ( .A(\b/SBOX[2].sbox/t[37] ), .B(\b/SBOX[2].sbox/y[3] ), .Z(
        \b/SBOX[2].sbox/z[10] ) );
  AND U2602 ( .A(\b/SBOX[2].sbox/t[44] ), .B(\b/SBOX[2].sbox/y[15] ), .Z(
        \b/SBOX[2].sbox/z[0] ) );
  AND U2603 ( .A(\b/SBOX[2].sbox/y[5] ), .B(\b/SBOX[2].sbox/y[1] ), .Z(
        \b/SBOX[2].sbox/t[8] ) );
  ANDN U2604 ( .A(\b/SBOX[2].sbox/y[16] ), .B(n1762), .Z(\b/SBOX[2].sbox/t[7] ) );
  XNOR U2605 ( .A(msg[17]), .B(msg[23]), .Z(n1762) );
  AND U2606 ( .A(\b/SBOX[2].sbox/y[4] ), .B(msg[16]), .Z(\b/SBOX[2].sbox/t[5] ) );
  AND U2607 ( .A(\b/SBOX[2].sbox/y[3] ), .B(\b/SBOX[2].sbox/y[6] ), .Z(
        \b/SBOX[2].sbox/t[3] ) );
  AND U2608 ( .A(\b/SBOX[2].sbox/t[38] ), .B(\b/SBOX[2].sbox/t[29] ), .Z(
        \b/SBOX[2].sbox/t[39] ) );
  AND U2609 ( .A(\b/SBOX[2].sbox/t[24] ), .B(n1763), .Z(\b/SBOX[2].sbox/t[36] ) );
  XOR U2610 ( .A(\b/SBOX[2].sbox/t[32] ), .B(\b/SBOX[2].sbox/t[26] ), .Z(n1763) );
  AND U2611 ( .A(\b/SBOX[2].sbox/t[31] ), .B(\b/SBOX[2].sbox/t[30] ), .Z(
        \b/SBOX[2].sbox/t[32] ) );
  AND U2612 ( .A(\b/SBOX[2].sbox/y[15] ), .B(\b/SBOX[2].sbox/y[12] ), .Z(
        \b/SBOX[2].sbox/t[2] ) );
  AND U2613 ( .A(\b/SBOX[2].sbox/t[27] ), .B(\b/SBOX[2].sbox/t[25] ), .Z(
        \b/SBOX[2].sbox/t[28] ) );
  AND U2614 ( .A(\b/SBOX[2].sbox/t[23] ), .B(\b/SBOX[2].sbox/t[21] ), .Z(
        \b/SBOX[2].sbox/t[26] ) );
  ANDN U2615 ( .A(\b/SBOX[2].sbox/y[10] ), .B(n1759), .Z(
        \b/SBOX[2].sbox/t[15] ) );
  XNOR U2616 ( .A(msg[18]), .B(msg[23]), .Z(n1759) );
  ANDN U2617 ( .A(\b/SBOX[2].sbox/y[17] ), .B(n1760), .Z(
        \b/SBOX[2].sbox/t[13] ) );
  XNOR U2618 ( .A(msg[18]), .B(msg[20]), .Z(n1760) );
  ANDN U2619 ( .A(\b/SBOX[2].sbox/y[11] ), .B(n1761), .Z(
        \b/SBOX[2].sbox/t[12] ) );
  XNOR U2620 ( .A(msg[20]), .B(msg[23]), .Z(n1761) );
  AND U2621 ( .A(\b/SBOX[2].sbox/y[2] ), .B(\b/SBOX[2].sbox/y[7] ), .Z(
        \b/SBOX[2].sbox/t[10] ) );
  AND U2622 ( .A(\b/SBOX[1].sbox/t[44] ), .B(\b/SBOX[1].sbox/y[12] ), .Z(
        \b/SBOX[1].sbox/z[9] ) );
  AND U2623 ( .A(\b/SBOX[1].sbox/t[41] ), .B(\b/SBOX[1].sbox/y[10] ), .Z(
        \b/SBOX[1].sbox/z[8] ) );
  AND U2624 ( .A(\b/SBOX[1].sbox/t[45] ), .B(\b/SBOX[1].sbox/y[17] ), .Z(
        \b/SBOX[1].sbox/z[7] ) );
  AND U2625 ( .A(\b/SBOX[1].sbox/t[42] ), .B(\b/SBOX[1].sbox/y[11] ), .Z(
        \b/SBOX[1].sbox/z[6] ) );
  AND U2626 ( .A(\b/SBOX[1].sbox/t[29] ), .B(\b/SBOX[1].sbox/y[7] ), .Z(
        \b/SBOX[1].sbox/z[5] ) );
  AND U2627 ( .A(\b/SBOX[1].sbox/t[40] ), .B(\b/SBOX[1].sbox/y[1] ), .Z(
        \b/SBOX[1].sbox/z[4] ) );
  AND U2628 ( .A(\b/SBOX[1].sbox/t[43] ), .B(\b/SBOX[1].sbox/y[16] ), .Z(
        \b/SBOX[1].sbox/z[3] ) );
  AND U2629 ( .A(msg[8]), .B(\b/SBOX[1].sbox/t[33] ), .Z(\b/SBOX[1].sbox/z[2] ) );
  AND U2630 ( .A(\b/SBOX[1].sbox/t[37] ), .B(\b/SBOX[1].sbox/y[6] ), .Z(
        \b/SBOX[1].sbox/z[1] ) );
  ANDN U2631 ( .A(\b/SBOX[1].sbox/t[41] ), .B(n1764), .Z(
        \b/SBOX[1].sbox/z[17] ) );
  ANDN U2632 ( .A(\b/SBOX[1].sbox/t[45] ), .B(n1765), .Z(
        \b/SBOX[1].sbox/z[16] ) );
  ANDN U2633 ( .A(\b/SBOX[1].sbox/t[42] ), .B(n1766), .Z(
        \b/SBOX[1].sbox/z[15] ) );
  AND U2634 ( .A(\b/SBOX[1].sbox/t[29] ), .B(\b/SBOX[1].sbox/y[2] ), .Z(
        \b/SBOX[1].sbox/z[14] ) );
  AND U2635 ( .A(\b/SBOX[1].sbox/t[40] ), .B(\b/SBOX[1].sbox/y[5] ), .Z(
        \b/SBOX[1].sbox/z[13] ) );
  ANDN U2636 ( .A(\b/SBOX[1].sbox/t[43] ), .B(n1767), .Z(
        \b/SBOX[1].sbox/z[12] ) );
  AND U2637 ( .A(\b/SBOX[1].sbox/t[33] ), .B(\b/SBOX[1].sbox/y[4] ), .Z(
        \b/SBOX[1].sbox/z[11] ) );
  AND U2638 ( .A(\b/SBOX[1].sbox/t[37] ), .B(\b/SBOX[1].sbox/y[3] ), .Z(
        \b/SBOX[1].sbox/z[10] ) );
  AND U2639 ( .A(\b/SBOX[1].sbox/t[44] ), .B(\b/SBOX[1].sbox/y[15] ), .Z(
        \b/SBOX[1].sbox/z[0] ) );
  AND U2640 ( .A(\b/SBOX[1].sbox/y[5] ), .B(\b/SBOX[1].sbox/y[1] ), .Z(
        \b/SBOX[1].sbox/t[8] ) );
  ANDN U2641 ( .A(\b/SBOX[1].sbox/y[16] ), .B(n1767), .Z(\b/SBOX[1].sbox/t[7] ) );
  XNOR U2642 ( .A(msg[15]), .B(msg[9]), .Z(n1767) );
  AND U2643 ( .A(\b/SBOX[1].sbox/y[4] ), .B(msg[8]), .Z(\b/SBOX[1].sbox/t[5] )
         );
  AND U2644 ( .A(\b/SBOX[1].sbox/y[3] ), .B(\b/SBOX[1].sbox/y[6] ), .Z(
        \b/SBOX[1].sbox/t[3] ) );
  AND U2645 ( .A(\b/SBOX[1].sbox/t[38] ), .B(\b/SBOX[1].sbox/t[29] ), .Z(
        \b/SBOX[1].sbox/t[39] ) );
  AND U2646 ( .A(\b/SBOX[1].sbox/t[24] ), .B(n1768), .Z(\b/SBOX[1].sbox/t[36] ) );
  XOR U2647 ( .A(\b/SBOX[1].sbox/t[32] ), .B(\b/SBOX[1].sbox/t[26] ), .Z(n1768) );
  AND U2648 ( .A(\b/SBOX[1].sbox/t[31] ), .B(\b/SBOX[1].sbox/t[30] ), .Z(
        \b/SBOX[1].sbox/t[32] ) );
  AND U2649 ( .A(\b/SBOX[1].sbox/y[15] ), .B(\b/SBOX[1].sbox/y[12] ), .Z(
        \b/SBOX[1].sbox/t[2] ) );
  AND U2650 ( .A(\b/SBOX[1].sbox/t[27] ), .B(\b/SBOX[1].sbox/t[25] ), .Z(
        \b/SBOX[1].sbox/t[28] ) );
  AND U2651 ( .A(\b/SBOX[1].sbox/t[23] ), .B(\b/SBOX[1].sbox/t[21] ), .Z(
        \b/SBOX[1].sbox/t[26] ) );
  ANDN U2652 ( .A(\b/SBOX[1].sbox/y[10] ), .B(n1764), .Z(
        \b/SBOX[1].sbox/t[15] ) );
  XNOR U2653 ( .A(msg[10]), .B(msg[15]), .Z(n1764) );
  ANDN U2654 ( .A(\b/SBOX[1].sbox/y[17] ), .B(n1765), .Z(
        \b/SBOX[1].sbox/t[13] ) );
  XNOR U2655 ( .A(msg[10]), .B(msg[12]), .Z(n1765) );
  ANDN U2656 ( .A(\b/SBOX[1].sbox/y[11] ), .B(n1766), .Z(
        \b/SBOX[1].sbox/t[12] ) );
  XNOR U2657 ( .A(msg[12]), .B(msg[15]), .Z(n1766) );
  AND U2658 ( .A(\b/SBOX[1].sbox/y[2] ), .B(\b/SBOX[1].sbox/y[7] ), .Z(
        \b/SBOX[1].sbox/t[10] ) );
  AND U2659 ( .A(\b/SBOX[15].sbox/t[44] ), .B(\b/SBOX[15].sbox/y[12] ), .Z(
        \b/SBOX[15].sbox/z[9] ) );
  AND U2660 ( .A(\b/SBOX[15].sbox/t[41] ), .B(\b/SBOX[15].sbox/y[10] ), .Z(
        \b/SBOX[15].sbox/z[8] ) );
  AND U2661 ( .A(\b/SBOX[15].sbox/t[45] ), .B(\b/SBOX[15].sbox/y[17] ), .Z(
        \b/SBOX[15].sbox/z[7] ) );
  AND U2662 ( .A(\b/SBOX[15].sbox/t[42] ), .B(\b/SBOX[15].sbox/y[11] ), .Z(
        \b/SBOX[15].sbox/z[6] ) );
  AND U2663 ( .A(\b/SBOX[15].sbox/t[29] ), .B(\b/SBOX[15].sbox/y[7] ), .Z(
        \b/SBOX[15].sbox/z[5] ) );
  AND U2664 ( .A(\b/SBOX[15].sbox/t[40] ), .B(\b/SBOX[15].sbox/y[1] ), .Z(
        \b/SBOX[15].sbox/z[4] ) );
  AND U2665 ( .A(\b/SBOX[15].sbox/t[43] ), .B(\b/SBOX[15].sbox/y[16] ), .Z(
        \b/SBOX[15].sbox/z[3] ) );
  AND U2666 ( .A(msg[120]), .B(\b/SBOX[15].sbox/t[33] ), .Z(
        \b/SBOX[15].sbox/z[2] ) );
  AND U2667 ( .A(\b/SBOX[15].sbox/t[37] ), .B(\b/SBOX[15].sbox/y[6] ), .Z(
        \b/SBOX[15].sbox/z[1] ) );
  ANDN U2668 ( .A(\b/SBOX[15].sbox/t[41] ), .B(n1769), .Z(
        \b/SBOX[15].sbox/z[17] ) );
  ANDN U2669 ( .A(\b/SBOX[15].sbox/t[45] ), .B(n1770), .Z(
        \b/SBOX[15].sbox/z[16] ) );
  ANDN U2670 ( .A(\b/SBOX[15].sbox/t[42] ), .B(n1771), .Z(
        \b/SBOX[15].sbox/z[15] ) );
  AND U2671 ( .A(\b/SBOX[15].sbox/t[29] ), .B(\b/SBOX[15].sbox/y[2] ), .Z(
        \b/SBOX[15].sbox/z[14] ) );
  AND U2672 ( .A(\b/SBOX[15].sbox/t[40] ), .B(\b/SBOX[15].sbox/y[5] ), .Z(
        \b/SBOX[15].sbox/z[13] ) );
  ANDN U2673 ( .A(\b/SBOX[15].sbox/t[43] ), .B(n1772), .Z(
        \b/SBOX[15].sbox/z[12] ) );
  AND U2674 ( .A(\b/SBOX[15].sbox/t[33] ), .B(\b/SBOX[15].sbox/y[4] ), .Z(
        \b/SBOX[15].sbox/z[11] ) );
  AND U2675 ( .A(\b/SBOX[15].sbox/t[37] ), .B(\b/SBOX[15].sbox/y[3] ), .Z(
        \b/SBOX[15].sbox/z[10] ) );
  AND U2676 ( .A(\b/SBOX[15].sbox/t[44] ), .B(\b/SBOX[15].sbox/y[15] ), .Z(
        \b/SBOX[15].sbox/z[0] ) );
  AND U2677 ( .A(\b/SBOX[15].sbox/y[5] ), .B(\b/SBOX[15].sbox/y[1] ), .Z(
        \b/SBOX[15].sbox/t[8] ) );
  ANDN U2678 ( .A(\b/SBOX[15].sbox/y[16] ), .B(n1772), .Z(
        \b/SBOX[15].sbox/t[7] ) );
  XNOR U2679 ( .A(msg[121]), .B(msg[127]), .Z(n1772) );
  AND U2680 ( .A(\b/SBOX[15].sbox/y[4] ), .B(msg[120]), .Z(
        \b/SBOX[15].sbox/t[5] ) );
  AND U2681 ( .A(\b/SBOX[15].sbox/y[3] ), .B(\b/SBOX[15].sbox/y[6] ), .Z(
        \b/SBOX[15].sbox/t[3] ) );
  AND U2682 ( .A(\b/SBOX[15].sbox/t[38] ), .B(\b/SBOX[15].sbox/t[29] ), .Z(
        \b/SBOX[15].sbox/t[39] ) );
  AND U2683 ( .A(\b/SBOX[15].sbox/t[24] ), .B(n1773), .Z(
        \b/SBOX[15].sbox/t[36] ) );
  XOR U2684 ( .A(\b/SBOX[15].sbox/t[32] ), .B(\b/SBOX[15].sbox/t[26] ), .Z(
        n1773) );
  AND U2685 ( .A(\b/SBOX[15].sbox/t[31] ), .B(\b/SBOX[15].sbox/t[30] ), .Z(
        \b/SBOX[15].sbox/t[32] ) );
  AND U2686 ( .A(\b/SBOX[15].sbox/y[15] ), .B(\b/SBOX[15].sbox/y[12] ), .Z(
        \b/SBOX[15].sbox/t[2] ) );
  AND U2687 ( .A(\b/SBOX[15].sbox/t[27] ), .B(\b/SBOX[15].sbox/t[25] ), .Z(
        \b/SBOX[15].sbox/t[28] ) );
  AND U2688 ( .A(\b/SBOX[15].sbox/t[23] ), .B(\b/SBOX[15].sbox/t[21] ), .Z(
        \b/SBOX[15].sbox/t[26] ) );
  ANDN U2689 ( .A(\b/SBOX[15].sbox/y[10] ), .B(n1769), .Z(
        \b/SBOX[15].sbox/t[15] ) );
  XNOR U2690 ( .A(msg[122]), .B(msg[127]), .Z(n1769) );
  ANDN U2691 ( .A(\b/SBOX[15].sbox/y[17] ), .B(n1770), .Z(
        \b/SBOX[15].sbox/t[13] ) );
  XNOR U2692 ( .A(msg[122]), .B(msg[124]), .Z(n1770) );
  ANDN U2693 ( .A(\b/SBOX[15].sbox/y[11] ), .B(n1771), .Z(
        \b/SBOX[15].sbox/t[12] ) );
  XNOR U2694 ( .A(msg[124]), .B(msg[127]), .Z(n1771) );
  AND U2695 ( .A(\b/SBOX[15].sbox/y[2] ), .B(\b/SBOX[15].sbox/y[7] ), .Z(
        \b/SBOX[15].sbox/t[10] ) );
  AND U2696 ( .A(\b/SBOX[14].sbox/t[44] ), .B(\b/SBOX[14].sbox/y[12] ), .Z(
        \b/SBOX[14].sbox/z[9] ) );
  AND U2697 ( .A(\b/SBOX[14].sbox/t[41] ), .B(\b/SBOX[14].sbox/y[10] ), .Z(
        \b/SBOX[14].sbox/z[8] ) );
  AND U2698 ( .A(\b/SBOX[14].sbox/t[45] ), .B(\b/SBOX[14].sbox/y[17] ), .Z(
        \b/SBOX[14].sbox/z[7] ) );
  AND U2699 ( .A(\b/SBOX[14].sbox/t[42] ), .B(\b/SBOX[14].sbox/y[11] ), .Z(
        \b/SBOX[14].sbox/z[6] ) );
  AND U2700 ( .A(\b/SBOX[14].sbox/t[29] ), .B(\b/SBOX[14].sbox/y[7] ), .Z(
        \b/SBOX[14].sbox/z[5] ) );
  AND U2701 ( .A(\b/SBOX[14].sbox/t[40] ), .B(\b/SBOX[14].sbox/y[1] ), .Z(
        \b/SBOX[14].sbox/z[4] ) );
  AND U2702 ( .A(\b/SBOX[14].sbox/t[43] ), .B(\b/SBOX[14].sbox/y[16] ), .Z(
        \b/SBOX[14].sbox/z[3] ) );
  AND U2703 ( .A(msg[112]), .B(\b/SBOX[14].sbox/t[33] ), .Z(
        \b/SBOX[14].sbox/z[2] ) );
  AND U2704 ( .A(\b/SBOX[14].sbox/t[37] ), .B(\b/SBOX[14].sbox/y[6] ), .Z(
        \b/SBOX[14].sbox/z[1] ) );
  ANDN U2705 ( .A(\b/SBOX[14].sbox/t[41] ), .B(n1774), .Z(
        \b/SBOX[14].sbox/z[17] ) );
  ANDN U2706 ( .A(\b/SBOX[14].sbox/t[45] ), .B(n1775), .Z(
        \b/SBOX[14].sbox/z[16] ) );
  ANDN U2707 ( .A(\b/SBOX[14].sbox/t[42] ), .B(n1776), .Z(
        \b/SBOX[14].sbox/z[15] ) );
  AND U2708 ( .A(\b/SBOX[14].sbox/t[29] ), .B(\b/SBOX[14].sbox/y[2] ), .Z(
        \b/SBOX[14].sbox/z[14] ) );
  AND U2709 ( .A(\b/SBOX[14].sbox/t[40] ), .B(\b/SBOX[14].sbox/y[5] ), .Z(
        \b/SBOX[14].sbox/z[13] ) );
  ANDN U2710 ( .A(\b/SBOX[14].sbox/t[43] ), .B(n1777), .Z(
        \b/SBOX[14].sbox/z[12] ) );
  AND U2711 ( .A(\b/SBOX[14].sbox/t[33] ), .B(\b/SBOX[14].sbox/y[4] ), .Z(
        \b/SBOX[14].sbox/z[11] ) );
  AND U2712 ( .A(\b/SBOX[14].sbox/t[37] ), .B(\b/SBOX[14].sbox/y[3] ), .Z(
        \b/SBOX[14].sbox/z[10] ) );
  AND U2713 ( .A(\b/SBOX[14].sbox/t[44] ), .B(\b/SBOX[14].sbox/y[15] ), .Z(
        \b/SBOX[14].sbox/z[0] ) );
  AND U2714 ( .A(\b/SBOX[14].sbox/y[5] ), .B(\b/SBOX[14].sbox/y[1] ), .Z(
        \b/SBOX[14].sbox/t[8] ) );
  ANDN U2715 ( .A(\b/SBOX[14].sbox/y[16] ), .B(n1777), .Z(
        \b/SBOX[14].sbox/t[7] ) );
  XNOR U2716 ( .A(msg[113]), .B(msg[119]), .Z(n1777) );
  AND U2717 ( .A(\b/SBOX[14].sbox/y[4] ), .B(msg[112]), .Z(
        \b/SBOX[14].sbox/t[5] ) );
  AND U2718 ( .A(\b/SBOX[14].sbox/y[3] ), .B(\b/SBOX[14].sbox/y[6] ), .Z(
        \b/SBOX[14].sbox/t[3] ) );
  AND U2719 ( .A(\b/SBOX[14].sbox/t[38] ), .B(\b/SBOX[14].sbox/t[29] ), .Z(
        \b/SBOX[14].sbox/t[39] ) );
  AND U2720 ( .A(\b/SBOX[14].sbox/t[24] ), .B(n1778), .Z(
        \b/SBOX[14].sbox/t[36] ) );
  XOR U2721 ( .A(\b/SBOX[14].sbox/t[32] ), .B(\b/SBOX[14].sbox/t[26] ), .Z(
        n1778) );
  AND U2722 ( .A(\b/SBOX[14].sbox/t[31] ), .B(\b/SBOX[14].sbox/t[30] ), .Z(
        \b/SBOX[14].sbox/t[32] ) );
  AND U2723 ( .A(\b/SBOX[14].sbox/y[15] ), .B(\b/SBOX[14].sbox/y[12] ), .Z(
        \b/SBOX[14].sbox/t[2] ) );
  AND U2724 ( .A(\b/SBOX[14].sbox/t[27] ), .B(\b/SBOX[14].sbox/t[25] ), .Z(
        \b/SBOX[14].sbox/t[28] ) );
  AND U2725 ( .A(\b/SBOX[14].sbox/t[23] ), .B(\b/SBOX[14].sbox/t[21] ), .Z(
        \b/SBOX[14].sbox/t[26] ) );
  ANDN U2726 ( .A(\b/SBOX[14].sbox/y[10] ), .B(n1774), .Z(
        \b/SBOX[14].sbox/t[15] ) );
  XNOR U2727 ( .A(msg[114]), .B(msg[119]), .Z(n1774) );
  ANDN U2728 ( .A(\b/SBOX[14].sbox/y[17] ), .B(n1775), .Z(
        \b/SBOX[14].sbox/t[13] ) );
  XNOR U2729 ( .A(msg[114]), .B(msg[116]), .Z(n1775) );
  ANDN U2730 ( .A(\b/SBOX[14].sbox/y[11] ), .B(n1776), .Z(
        \b/SBOX[14].sbox/t[12] ) );
  XNOR U2731 ( .A(msg[116]), .B(msg[119]), .Z(n1776) );
  AND U2732 ( .A(\b/SBOX[14].sbox/y[2] ), .B(\b/SBOX[14].sbox/y[7] ), .Z(
        \b/SBOX[14].sbox/t[10] ) );
  AND U2733 ( .A(\b/SBOX[13].sbox/t[44] ), .B(\b/SBOX[13].sbox/y[12] ), .Z(
        \b/SBOX[13].sbox/z[9] ) );
  AND U2734 ( .A(\b/SBOX[13].sbox/t[41] ), .B(\b/SBOX[13].sbox/y[10] ), .Z(
        \b/SBOX[13].sbox/z[8] ) );
  AND U2735 ( .A(\b/SBOX[13].sbox/t[45] ), .B(\b/SBOX[13].sbox/y[17] ), .Z(
        \b/SBOX[13].sbox/z[7] ) );
  AND U2736 ( .A(\b/SBOX[13].sbox/t[42] ), .B(\b/SBOX[13].sbox/y[11] ), .Z(
        \b/SBOX[13].sbox/z[6] ) );
  AND U2737 ( .A(\b/SBOX[13].sbox/t[29] ), .B(\b/SBOX[13].sbox/y[7] ), .Z(
        \b/SBOX[13].sbox/z[5] ) );
  AND U2738 ( .A(\b/SBOX[13].sbox/t[40] ), .B(\b/SBOX[13].sbox/y[1] ), .Z(
        \b/SBOX[13].sbox/z[4] ) );
  AND U2739 ( .A(\b/SBOX[13].sbox/t[43] ), .B(\b/SBOX[13].sbox/y[16] ), .Z(
        \b/SBOX[13].sbox/z[3] ) );
  AND U2740 ( .A(msg[104]), .B(\b/SBOX[13].sbox/t[33] ), .Z(
        \b/SBOX[13].sbox/z[2] ) );
  AND U2741 ( .A(\b/SBOX[13].sbox/t[37] ), .B(\b/SBOX[13].sbox/y[6] ), .Z(
        \b/SBOX[13].sbox/z[1] ) );
  ANDN U2742 ( .A(\b/SBOX[13].sbox/t[41] ), .B(n1779), .Z(
        \b/SBOX[13].sbox/z[17] ) );
  ANDN U2743 ( .A(\b/SBOX[13].sbox/t[45] ), .B(n1780), .Z(
        \b/SBOX[13].sbox/z[16] ) );
  ANDN U2744 ( .A(\b/SBOX[13].sbox/t[42] ), .B(n1781), .Z(
        \b/SBOX[13].sbox/z[15] ) );
  AND U2745 ( .A(\b/SBOX[13].sbox/t[29] ), .B(\b/SBOX[13].sbox/y[2] ), .Z(
        \b/SBOX[13].sbox/z[14] ) );
  AND U2746 ( .A(\b/SBOX[13].sbox/t[40] ), .B(\b/SBOX[13].sbox/y[5] ), .Z(
        \b/SBOX[13].sbox/z[13] ) );
  ANDN U2747 ( .A(\b/SBOX[13].sbox/t[43] ), .B(n1782), .Z(
        \b/SBOX[13].sbox/z[12] ) );
  AND U2748 ( .A(\b/SBOX[13].sbox/t[33] ), .B(\b/SBOX[13].sbox/y[4] ), .Z(
        \b/SBOX[13].sbox/z[11] ) );
  AND U2749 ( .A(\b/SBOX[13].sbox/t[37] ), .B(\b/SBOX[13].sbox/y[3] ), .Z(
        \b/SBOX[13].sbox/z[10] ) );
  AND U2750 ( .A(\b/SBOX[13].sbox/t[44] ), .B(\b/SBOX[13].sbox/y[15] ), .Z(
        \b/SBOX[13].sbox/z[0] ) );
  AND U2751 ( .A(\b/SBOX[13].sbox/y[5] ), .B(\b/SBOX[13].sbox/y[1] ), .Z(
        \b/SBOX[13].sbox/t[8] ) );
  ANDN U2752 ( .A(\b/SBOX[13].sbox/y[16] ), .B(n1782), .Z(
        \b/SBOX[13].sbox/t[7] ) );
  XNOR U2753 ( .A(msg[105]), .B(msg[111]), .Z(n1782) );
  AND U2754 ( .A(\b/SBOX[13].sbox/y[4] ), .B(msg[104]), .Z(
        \b/SBOX[13].sbox/t[5] ) );
  AND U2755 ( .A(\b/SBOX[13].sbox/y[3] ), .B(\b/SBOX[13].sbox/y[6] ), .Z(
        \b/SBOX[13].sbox/t[3] ) );
  AND U2756 ( .A(\b/SBOX[13].sbox/t[38] ), .B(\b/SBOX[13].sbox/t[29] ), .Z(
        \b/SBOX[13].sbox/t[39] ) );
  AND U2757 ( .A(\b/SBOX[13].sbox/t[24] ), .B(n1783), .Z(
        \b/SBOX[13].sbox/t[36] ) );
  XOR U2758 ( .A(\b/SBOX[13].sbox/t[32] ), .B(\b/SBOX[13].sbox/t[26] ), .Z(
        n1783) );
  AND U2759 ( .A(\b/SBOX[13].sbox/t[31] ), .B(\b/SBOX[13].sbox/t[30] ), .Z(
        \b/SBOX[13].sbox/t[32] ) );
  AND U2760 ( .A(\b/SBOX[13].sbox/y[15] ), .B(\b/SBOX[13].sbox/y[12] ), .Z(
        \b/SBOX[13].sbox/t[2] ) );
  AND U2761 ( .A(\b/SBOX[13].sbox/t[27] ), .B(\b/SBOX[13].sbox/t[25] ), .Z(
        \b/SBOX[13].sbox/t[28] ) );
  AND U2762 ( .A(\b/SBOX[13].sbox/t[23] ), .B(\b/SBOX[13].sbox/t[21] ), .Z(
        \b/SBOX[13].sbox/t[26] ) );
  ANDN U2763 ( .A(\b/SBOX[13].sbox/y[10] ), .B(n1779), .Z(
        \b/SBOX[13].sbox/t[15] ) );
  XNOR U2764 ( .A(msg[106]), .B(msg[111]), .Z(n1779) );
  ANDN U2765 ( .A(\b/SBOX[13].sbox/y[17] ), .B(n1780), .Z(
        \b/SBOX[13].sbox/t[13] ) );
  XNOR U2766 ( .A(msg[106]), .B(msg[108]), .Z(n1780) );
  ANDN U2767 ( .A(\b/SBOX[13].sbox/y[11] ), .B(n1781), .Z(
        \b/SBOX[13].sbox/t[12] ) );
  XNOR U2768 ( .A(msg[108]), .B(msg[111]), .Z(n1781) );
  AND U2769 ( .A(\b/SBOX[13].sbox/y[2] ), .B(\b/SBOX[13].sbox/y[7] ), .Z(
        \b/SBOX[13].sbox/t[10] ) );
  AND U2770 ( .A(\b/SBOX[12].sbox/t[44] ), .B(\b/SBOX[12].sbox/y[12] ), .Z(
        \b/SBOX[12].sbox/z[9] ) );
  AND U2771 ( .A(\b/SBOX[12].sbox/t[41] ), .B(\b/SBOX[12].sbox/y[10] ), .Z(
        \b/SBOX[12].sbox/z[8] ) );
  AND U2772 ( .A(\b/SBOX[12].sbox/t[45] ), .B(\b/SBOX[12].sbox/y[17] ), .Z(
        \b/SBOX[12].sbox/z[7] ) );
  AND U2773 ( .A(\b/SBOX[12].sbox/t[42] ), .B(\b/SBOX[12].sbox/y[11] ), .Z(
        \b/SBOX[12].sbox/z[6] ) );
  AND U2774 ( .A(\b/SBOX[12].sbox/t[29] ), .B(\b/SBOX[12].sbox/y[7] ), .Z(
        \b/SBOX[12].sbox/z[5] ) );
  AND U2775 ( .A(\b/SBOX[12].sbox/t[40] ), .B(\b/SBOX[12].sbox/y[1] ), .Z(
        \b/SBOX[12].sbox/z[4] ) );
  AND U2776 ( .A(\b/SBOX[12].sbox/t[43] ), .B(\b/SBOX[12].sbox/y[16] ), .Z(
        \b/SBOX[12].sbox/z[3] ) );
  AND U2777 ( .A(msg[96]), .B(\b/SBOX[12].sbox/t[33] ), .Z(
        \b/SBOX[12].sbox/z[2] ) );
  AND U2778 ( .A(\b/SBOX[12].sbox/t[37] ), .B(\b/SBOX[12].sbox/y[6] ), .Z(
        \b/SBOX[12].sbox/z[1] ) );
  ANDN U2779 ( .A(\b/SBOX[12].sbox/t[41] ), .B(n1784), .Z(
        \b/SBOX[12].sbox/z[17] ) );
  ANDN U2780 ( .A(\b/SBOX[12].sbox/t[45] ), .B(n1785), .Z(
        \b/SBOX[12].sbox/z[16] ) );
  ANDN U2781 ( .A(\b/SBOX[12].sbox/t[42] ), .B(n1786), .Z(
        \b/SBOX[12].sbox/z[15] ) );
  AND U2782 ( .A(\b/SBOX[12].sbox/t[29] ), .B(\b/SBOX[12].sbox/y[2] ), .Z(
        \b/SBOX[12].sbox/z[14] ) );
  AND U2783 ( .A(\b/SBOX[12].sbox/t[40] ), .B(\b/SBOX[12].sbox/y[5] ), .Z(
        \b/SBOX[12].sbox/z[13] ) );
  ANDN U2784 ( .A(\b/SBOX[12].sbox/t[43] ), .B(n1787), .Z(
        \b/SBOX[12].sbox/z[12] ) );
  AND U2785 ( .A(\b/SBOX[12].sbox/t[33] ), .B(\b/SBOX[12].sbox/y[4] ), .Z(
        \b/SBOX[12].sbox/z[11] ) );
  AND U2786 ( .A(\b/SBOX[12].sbox/t[37] ), .B(\b/SBOX[12].sbox/y[3] ), .Z(
        \b/SBOX[12].sbox/z[10] ) );
  AND U2787 ( .A(\b/SBOX[12].sbox/t[44] ), .B(\b/SBOX[12].sbox/y[15] ), .Z(
        \b/SBOX[12].sbox/z[0] ) );
  AND U2788 ( .A(\b/SBOX[12].sbox/y[5] ), .B(\b/SBOX[12].sbox/y[1] ), .Z(
        \b/SBOX[12].sbox/t[8] ) );
  ANDN U2789 ( .A(\b/SBOX[12].sbox/y[16] ), .B(n1787), .Z(
        \b/SBOX[12].sbox/t[7] ) );
  XNOR U2790 ( .A(msg[103]), .B(msg[97]), .Z(n1787) );
  AND U2791 ( .A(\b/SBOX[12].sbox/y[4] ), .B(msg[96]), .Z(
        \b/SBOX[12].sbox/t[5] ) );
  AND U2792 ( .A(\b/SBOX[12].sbox/y[3] ), .B(\b/SBOX[12].sbox/y[6] ), .Z(
        \b/SBOX[12].sbox/t[3] ) );
  AND U2793 ( .A(\b/SBOX[12].sbox/t[38] ), .B(\b/SBOX[12].sbox/t[29] ), .Z(
        \b/SBOX[12].sbox/t[39] ) );
  AND U2794 ( .A(\b/SBOX[12].sbox/t[24] ), .B(n1788), .Z(
        \b/SBOX[12].sbox/t[36] ) );
  XOR U2795 ( .A(\b/SBOX[12].sbox/t[32] ), .B(\b/SBOX[12].sbox/t[26] ), .Z(
        n1788) );
  AND U2796 ( .A(\b/SBOX[12].sbox/t[31] ), .B(\b/SBOX[12].sbox/t[30] ), .Z(
        \b/SBOX[12].sbox/t[32] ) );
  AND U2797 ( .A(\b/SBOX[12].sbox/y[15] ), .B(\b/SBOX[12].sbox/y[12] ), .Z(
        \b/SBOX[12].sbox/t[2] ) );
  AND U2798 ( .A(\b/SBOX[12].sbox/t[27] ), .B(\b/SBOX[12].sbox/t[25] ), .Z(
        \b/SBOX[12].sbox/t[28] ) );
  AND U2799 ( .A(\b/SBOX[12].sbox/t[23] ), .B(\b/SBOX[12].sbox/t[21] ), .Z(
        \b/SBOX[12].sbox/t[26] ) );
  ANDN U2800 ( .A(\b/SBOX[12].sbox/y[10] ), .B(n1784), .Z(
        \b/SBOX[12].sbox/t[15] ) );
  XNOR U2801 ( .A(msg[103]), .B(msg[98]), .Z(n1784) );
  ANDN U2802 ( .A(\b/SBOX[12].sbox/y[17] ), .B(n1785), .Z(
        \b/SBOX[12].sbox/t[13] ) );
  XNOR U2803 ( .A(msg[100]), .B(msg[98]), .Z(n1785) );
  ANDN U2804 ( .A(\b/SBOX[12].sbox/y[11] ), .B(n1786), .Z(
        \b/SBOX[12].sbox/t[12] ) );
  XNOR U2805 ( .A(msg[100]), .B(msg[103]), .Z(n1786) );
  AND U2806 ( .A(\b/SBOX[12].sbox/y[2] ), .B(\b/SBOX[12].sbox/y[7] ), .Z(
        \b/SBOX[12].sbox/t[10] ) );
  AND U2807 ( .A(\b/SBOX[11].sbox/t[44] ), .B(\b/SBOX[11].sbox/y[12] ), .Z(
        \b/SBOX[11].sbox/z[9] ) );
  AND U2808 ( .A(\b/SBOX[11].sbox/t[41] ), .B(\b/SBOX[11].sbox/y[10] ), .Z(
        \b/SBOX[11].sbox/z[8] ) );
  AND U2809 ( .A(\b/SBOX[11].sbox/t[45] ), .B(\b/SBOX[11].sbox/y[17] ), .Z(
        \b/SBOX[11].sbox/z[7] ) );
  AND U2810 ( .A(\b/SBOX[11].sbox/t[42] ), .B(\b/SBOX[11].sbox/y[11] ), .Z(
        \b/SBOX[11].sbox/z[6] ) );
  AND U2811 ( .A(\b/SBOX[11].sbox/t[29] ), .B(\b/SBOX[11].sbox/y[7] ), .Z(
        \b/SBOX[11].sbox/z[5] ) );
  AND U2812 ( .A(\b/SBOX[11].sbox/t[40] ), .B(\b/SBOX[11].sbox/y[1] ), .Z(
        \b/SBOX[11].sbox/z[4] ) );
  AND U2813 ( .A(\b/SBOX[11].sbox/t[43] ), .B(\b/SBOX[11].sbox/y[16] ), .Z(
        \b/SBOX[11].sbox/z[3] ) );
  AND U2814 ( .A(msg[88]), .B(\b/SBOX[11].sbox/t[33] ), .Z(
        \b/SBOX[11].sbox/z[2] ) );
  AND U2815 ( .A(\b/SBOX[11].sbox/t[37] ), .B(\b/SBOX[11].sbox/y[6] ), .Z(
        \b/SBOX[11].sbox/z[1] ) );
  ANDN U2816 ( .A(\b/SBOX[11].sbox/t[41] ), .B(n1789), .Z(
        \b/SBOX[11].sbox/z[17] ) );
  ANDN U2817 ( .A(\b/SBOX[11].sbox/t[45] ), .B(n1790), .Z(
        \b/SBOX[11].sbox/z[16] ) );
  ANDN U2818 ( .A(\b/SBOX[11].sbox/t[42] ), .B(n1791), .Z(
        \b/SBOX[11].sbox/z[15] ) );
  AND U2819 ( .A(\b/SBOX[11].sbox/t[29] ), .B(\b/SBOX[11].sbox/y[2] ), .Z(
        \b/SBOX[11].sbox/z[14] ) );
  AND U2820 ( .A(\b/SBOX[11].sbox/t[40] ), .B(\b/SBOX[11].sbox/y[5] ), .Z(
        \b/SBOX[11].sbox/z[13] ) );
  ANDN U2821 ( .A(\b/SBOX[11].sbox/t[43] ), .B(n1792), .Z(
        \b/SBOX[11].sbox/z[12] ) );
  AND U2822 ( .A(\b/SBOX[11].sbox/t[33] ), .B(\b/SBOX[11].sbox/y[4] ), .Z(
        \b/SBOX[11].sbox/z[11] ) );
  AND U2823 ( .A(\b/SBOX[11].sbox/t[37] ), .B(\b/SBOX[11].sbox/y[3] ), .Z(
        \b/SBOX[11].sbox/z[10] ) );
  AND U2824 ( .A(\b/SBOX[11].sbox/t[44] ), .B(\b/SBOX[11].sbox/y[15] ), .Z(
        \b/SBOX[11].sbox/z[0] ) );
  AND U2825 ( .A(\b/SBOX[11].sbox/y[5] ), .B(\b/SBOX[11].sbox/y[1] ), .Z(
        \b/SBOX[11].sbox/t[8] ) );
  ANDN U2826 ( .A(\b/SBOX[11].sbox/y[16] ), .B(n1792), .Z(
        \b/SBOX[11].sbox/t[7] ) );
  XNOR U2827 ( .A(msg[89]), .B(msg[95]), .Z(n1792) );
  AND U2828 ( .A(\b/SBOX[11].sbox/y[4] ), .B(msg[88]), .Z(
        \b/SBOX[11].sbox/t[5] ) );
  AND U2829 ( .A(\b/SBOX[11].sbox/y[3] ), .B(\b/SBOX[11].sbox/y[6] ), .Z(
        \b/SBOX[11].sbox/t[3] ) );
  AND U2830 ( .A(\b/SBOX[11].sbox/t[38] ), .B(\b/SBOX[11].sbox/t[29] ), .Z(
        \b/SBOX[11].sbox/t[39] ) );
  AND U2831 ( .A(\b/SBOX[11].sbox/t[24] ), .B(n1793), .Z(
        \b/SBOX[11].sbox/t[36] ) );
  XOR U2832 ( .A(\b/SBOX[11].sbox/t[32] ), .B(\b/SBOX[11].sbox/t[26] ), .Z(
        n1793) );
  AND U2833 ( .A(\b/SBOX[11].sbox/t[31] ), .B(\b/SBOX[11].sbox/t[30] ), .Z(
        \b/SBOX[11].sbox/t[32] ) );
  AND U2834 ( .A(\b/SBOX[11].sbox/y[15] ), .B(\b/SBOX[11].sbox/y[12] ), .Z(
        \b/SBOX[11].sbox/t[2] ) );
  AND U2835 ( .A(\b/SBOX[11].sbox/t[27] ), .B(\b/SBOX[11].sbox/t[25] ), .Z(
        \b/SBOX[11].sbox/t[28] ) );
  AND U2836 ( .A(\b/SBOX[11].sbox/t[23] ), .B(\b/SBOX[11].sbox/t[21] ), .Z(
        \b/SBOX[11].sbox/t[26] ) );
  ANDN U2837 ( .A(\b/SBOX[11].sbox/y[10] ), .B(n1789), .Z(
        \b/SBOX[11].sbox/t[15] ) );
  XNOR U2838 ( .A(msg[90]), .B(msg[95]), .Z(n1789) );
  ANDN U2839 ( .A(\b/SBOX[11].sbox/y[17] ), .B(n1790), .Z(
        \b/SBOX[11].sbox/t[13] ) );
  XNOR U2840 ( .A(msg[90]), .B(msg[92]), .Z(n1790) );
  ANDN U2841 ( .A(\b/SBOX[11].sbox/y[11] ), .B(n1791), .Z(
        \b/SBOX[11].sbox/t[12] ) );
  XNOR U2842 ( .A(msg[92]), .B(msg[95]), .Z(n1791) );
  AND U2843 ( .A(\b/SBOX[11].sbox/y[2] ), .B(\b/SBOX[11].sbox/y[7] ), .Z(
        \b/SBOX[11].sbox/t[10] ) );
  AND U2844 ( .A(\b/SBOX[10].sbox/t[44] ), .B(\b/SBOX[10].sbox/y[12] ), .Z(
        \b/SBOX[10].sbox/z[9] ) );
  AND U2845 ( .A(\b/SBOX[10].sbox/t[41] ), .B(\b/SBOX[10].sbox/y[10] ), .Z(
        \b/SBOX[10].sbox/z[8] ) );
  AND U2846 ( .A(\b/SBOX[10].sbox/t[45] ), .B(\b/SBOX[10].sbox/y[17] ), .Z(
        \b/SBOX[10].sbox/z[7] ) );
  AND U2847 ( .A(\b/SBOX[10].sbox/t[42] ), .B(\b/SBOX[10].sbox/y[11] ), .Z(
        \b/SBOX[10].sbox/z[6] ) );
  AND U2848 ( .A(\b/SBOX[10].sbox/t[29] ), .B(\b/SBOX[10].sbox/y[7] ), .Z(
        \b/SBOX[10].sbox/z[5] ) );
  AND U2849 ( .A(\b/SBOX[10].sbox/t[40] ), .B(\b/SBOX[10].sbox/y[1] ), .Z(
        \b/SBOX[10].sbox/z[4] ) );
  AND U2850 ( .A(\b/SBOX[10].sbox/t[43] ), .B(\b/SBOX[10].sbox/y[16] ), .Z(
        \b/SBOX[10].sbox/z[3] ) );
  AND U2851 ( .A(msg[80]), .B(\b/SBOX[10].sbox/t[33] ), .Z(
        \b/SBOX[10].sbox/z[2] ) );
  AND U2852 ( .A(\b/SBOX[10].sbox/t[37] ), .B(\b/SBOX[10].sbox/y[6] ), .Z(
        \b/SBOX[10].sbox/z[1] ) );
  ANDN U2853 ( .A(\b/SBOX[10].sbox/t[41] ), .B(n1794), .Z(
        \b/SBOX[10].sbox/z[17] ) );
  ANDN U2854 ( .A(\b/SBOX[10].sbox/t[45] ), .B(n1795), .Z(
        \b/SBOX[10].sbox/z[16] ) );
  ANDN U2855 ( .A(\b/SBOX[10].sbox/t[42] ), .B(n1796), .Z(
        \b/SBOX[10].sbox/z[15] ) );
  AND U2856 ( .A(\b/SBOX[10].sbox/t[29] ), .B(\b/SBOX[10].sbox/y[2] ), .Z(
        \b/SBOX[10].sbox/z[14] ) );
  AND U2857 ( .A(\b/SBOX[10].sbox/t[40] ), .B(\b/SBOX[10].sbox/y[5] ), .Z(
        \b/SBOX[10].sbox/z[13] ) );
  ANDN U2858 ( .A(\b/SBOX[10].sbox/t[43] ), .B(n1797), .Z(
        \b/SBOX[10].sbox/z[12] ) );
  AND U2859 ( .A(\b/SBOX[10].sbox/t[33] ), .B(\b/SBOX[10].sbox/y[4] ), .Z(
        \b/SBOX[10].sbox/z[11] ) );
  AND U2860 ( .A(\b/SBOX[10].sbox/t[37] ), .B(\b/SBOX[10].sbox/y[3] ), .Z(
        \b/SBOX[10].sbox/z[10] ) );
  AND U2861 ( .A(\b/SBOX[10].sbox/t[44] ), .B(\b/SBOX[10].sbox/y[15] ), .Z(
        \b/SBOX[10].sbox/z[0] ) );
  AND U2862 ( .A(\b/SBOX[10].sbox/y[5] ), .B(\b/SBOX[10].sbox/y[1] ), .Z(
        \b/SBOX[10].sbox/t[8] ) );
  ANDN U2863 ( .A(\b/SBOX[10].sbox/y[16] ), .B(n1797), .Z(
        \b/SBOX[10].sbox/t[7] ) );
  XNOR U2864 ( .A(msg[81]), .B(msg[87]), .Z(n1797) );
  AND U2865 ( .A(\b/SBOX[10].sbox/y[4] ), .B(msg[80]), .Z(
        \b/SBOX[10].sbox/t[5] ) );
  AND U2866 ( .A(\b/SBOX[10].sbox/y[3] ), .B(\b/SBOX[10].sbox/y[6] ), .Z(
        \b/SBOX[10].sbox/t[3] ) );
  AND U2867 ( .A(\b/SBOX[10].sbox/t[38] ), .B(\b/SBOX[10].sbox/t[29] ), .Z(
        \b/SBOX[10].sbox/t[39] ) );
  AND U2868 ( .A(\b/SBOX[10].sbox/t[24] ), .B(n1798), .Z(
        \b/SBOX[10].sbox/t[36] ) );
  XOR U2869 ( .A(\b/SBOX[10].sbox/t[32] ), .B(\b/SBOX[10].sbox/t[26] ), .Z(
        n1798) );
  AND U2870 ( .A(\b/SBOX[10].sbox/t[31] ), .B(\b/SBOX[10].sbox/t[30] ), .Z(
        \b/SBOX[10].sbox/t[32] ) );
  AND U2871 ( .A(\b/SBOX[10].sbox/y[15] ), .B(\b/SBOX[10].sbox/y[12] ), .Z(
        \b/SBOX[10].sbox/t[2] ) );
  AND U2872 ( .A(\b/SBOX[10].sbox/t[27] ), .B(\b/SBOX[10].sbox/t[25] ), .Z(
        \b/SBOX[10].sbox/t[28] ) );
  AND U2873 ( .A(\b/SBOX[10].sbox/t[23] ), .B(\b/SBOX[10].sbox/t[21] ), .Z(
        \b/SBOX[10].sbox/t[26] ) );
  ANDN U2874 ( .A(\b/SBOX[10].sbox/y[10] ), .B(n1794), .Z(
        \b/SBOX[10].sbox/t[15] ) );
  XNOR U2875 ( .A(msg[82]), .B(msg[87]), .Z(n1794) );
  ANDN U2876 ( .A(\b/SBOX[10].sbox/y[17] ), .B(n1795), .Z(
        \b/SBOX[10].sbox/t[13] ) );
  XNOR U2877 ( .A(msg[82]), .B(msg[84]), .Z(n1795) );
  ANDN U2878 ( .A(\b/SBOX[10].sbox/y[11] ), .B(n1796), .Z(
        \b/SBOX[10].sbox/t[12] ) );
  XNOR U2879 ( .A(msg[84]), .B(msg[87]), .Z(n1796) );
  AND U2880 ( .A(\b/SBOX[10].sbox/y[2] ), .B(\b/SBOX[10].sbox/y[7] ), .Z(
        \b/SBOX[10].sbox/t[10] ) );
  AND U2881 ( .A(\b/SBOX[0].sbox/t[44] ), .B(\b/SBOX[0].sbox/y[12] ), .Z(
        \b/SBOX[0].sbox/z[9] ) );
  AND U2882 ( .A(\b/SBOX[0].sbox/t[41] ), .B(\b/SBOX[0].sbox/y[10] ), .Z(
        \b/SBOX[0].sbox/z[8] ) );
  AND U2883 ( .A(\b/SBOX[0].sbox/t[45] ), .B(\b/SBOX[0].sbox/y[17] ), .Z(
        \b/SBOX[0].sbox/z[7] ) );
  AND U2884 ( .A(\b/SBOX[0].sbox/t[42] ), .B(\b/SBOX[0].sbox/y[11] ), .Z(
        \b/SBOX[0].sbox/z[6] ) );
  AND U2885 ( .A(\b/SBOX[0].sbox/t[29] ), .B(\b/SBOX[0].sbox/y[7] ), .Z(
        \b/SBOX[0].sbox/z[5] ) );
  AND U2886 ( .A(\b/SBOX[0].sbox/t[40] ), .B(\b/SBOX[0].sbox/y[1] ), .Z(
        \b/SBOX[0].sbox/z[4] ) );
  AND U2887 ( .A(\b/SBOX[0].sbox/t[43] ), .B(\b/SBOX[0].sbox/y[16] ), .Z(
        \b/SBOX[0].sbox/z[3] ) );
  AND U2888 ( .A(msg[0]), .B(\b/SBOX[0].sbox/t[33] ), .Z(\b/SBOX[0].sbox/z[2] ) );
  AND U2889 ( .A(\b/SBOX[0].sbox/t[37] ), .B(\b/SBOX[0].sbox/y[6] ), .Z(
        \b/SBOX[0].sbox/z[1] ) );
  ANDN U2890 ( .A(\b/SBOX[0].sbox/t[41] ), .B(n1799), .Z(
        \b/SBOX[0].sbox/z[17] ) );
  ANDN U2891 ( .A(\b/SBOX[0].sbox/t[45] ), .B(n1800), .Z(
        \b/SBOX[0].sbox/z[16] ) );
  ANDN U2892 ( .A(\b/SBOX[0].sbox/t[42] ), .B(n1801), .Z(
        \b/SBOX[0].sbox/z[15] ) );
  AND U2893 ( .A(\b/SBOX[0].sbox/t[29] ), .B(\b/SBOX[0].sbox/y[2] ), .Z(
        \b/SBOX[0].sbox/z[14] ) );
  AND U2894 ( .A(\b/SBOX[0].sbox/t[40] ), .B(\b/SBOX[0].sbox/y[5] ), .Z(
        \b/SBOX[0].sbox/z[13] ) );
  ANDN U2895 ( .A(\b/SBOX[0].sbox/t[43] ), .B(n1802), .Z(
        \b/SBOX[0].sbox/z[12] ) );
  AND U2896 ( .A(\b/SBOX[0].sbox/t[33] ), .B(\b/SBOX[0].sbox/y[4] ), .Z(
        \b/SBOX[0].sbox/z[11] ) );
  AND U2897 ( .A(\b/SBOX[0].sbox/t[37] ), .B(\b/SBOX[0].sbox/y[3] ), .Z(
        \b/SBOX[0].sbox/z[10] ) );
  AND U2898 ( .A(\b/SBOX[0].sbox/t[44] ), .B(\b/SBOX[0].sbox/y[15] ), .Z(
        \b/SBOX[0].sbox/z[0] ) );
  AND U2899 ( .A(\b/SBOX[0].sbox/y[5] ), .B(\b/SBOX[0].sbox/y[1] ), .Z(
        \b/SBOX[0].sbox/t[8] ) );
  ANDN U2900 ( .A(\b/SBOX[0].sbox/y[16] ), .B(n1802), .Z(\b/SBOX[0].sbox/t[7] ) );
  XNOR U2901 ( .A(msg[1]), .B(msg[7]), .Z(n1802) );
  AND U2902 ( .A(\b/SBOX[0].sbox/y[4] ), .B(msg[0]), .Z(\b/SBOX[0].sbox/t[5] )
         );
  AND U2903 ( .A(\b/SBOX[0].sbox/y[3] ), .B(\b/SBOX[0].sbox/y[6] ), .Z(
        \b/SBOX[0].sbox/t[3] ) );
  AND U2904 ( .A(\b/SBOX[0].sbox/t[38] ), .B(\b/SBOX[0].sbox/t[29] ), .Z(
        \b/SBOX[0].sbox/t[39] ) );
  AND U2905 ( .A(\b/SBOX[0].sbox/t[24] ), .B(n1803), .Z(\b/SBOX[0].sbox/t[36] ) );
  XOR U2906 ( .A(\b/SBOX[0].sbox/t[32] ), .B(\b/SBOX[0].sbox/t[26] ), .Z(n1803) );
  AND U2907 ( .A(\b/SBOX[0].sbox/t[31] ), .B(\b/SBOX[0].sbox/t[30] ), .Z(
        \b/SBOX[0].sbox/t[32] ) );
  AND U2908 ( .A(\b/SBOX[0].sbox/y[15] ), .B(\b/SBOX[0].sbox/y[12] ), .Z(
        \b/SBOX[0].sbox/t[2] ) );
  AND U2909 ( .A(\b/SBOX[0].sbox/t[27] ), .B(\b/SBOX[0].sbox/t[25] ), .Z(
        \b/SBOX[0].sbox/t[28] ) );
  AND U2910 ( .A(\b/SBOX[0].sbox/t[23] ), .B(\b/SBOX[0].sbox/t[21] ), .Z(
        \b/SBOX[0].sbox/t[26] ) );
  ANDN U2911 ( .A(\b/SBOX[0].sbox/y[10] ), .B(n1799), .Z(
        \b/SBOX[0].sbox/t[15] ) );
  XNOR U2912 ( .A(msg[2]), .B(msg[7]), .Z(n1799) );
  ANDN U2913 ( .A(\b/SBOX[0].sbox/y[17] ), .B(n1800), .Z(
        \b/SBOX[0].sbox/t[13] ) );
  XNOR U2914 ( .A(msg[2]), .B(msg[4]), .Z(n1800) );
  ANDN U2915 ( .A(\b/SBOX[0].sbox/y[11] ), .B(n1801), .Z(
        \b/SBOX[0].sbox/t[12] ) );
  XNOR U2916 ( .A(msg[4]), .B(msg[7]), .Z(n1801) );
  AND U2917 ( .A(\b/SBOX[0].sbox/y[2] ), .B(\b/SBOX[0].sbox/y[7] ), .Z(
        \b/SBOX[0].sbox/t[10] ) );
  XNOR U2918 ( .A(n1700), .B(n1804), .Z(N7) );
  NOR U2919 ( .A(n1685), .B(n1805), .Z(n1804) );
  IV U2920 ( .A(counter[2]), .Z(n1685) );
  IV U2921 ( .A(counter[3]), .Z(n1700) );
  XNOR U2922 ( .A(counter[2]), .B(n1805), .Z(N6) );
  NANDN U2923 ( .B(n1689), .A(counter[0]), .Z(n1805) );
  XNOR U2924 ( .A(n1689), .B(counter[0]), .Z(N5) );
  IV U2925 ( .A(counter[1]), .Z(n1689) );
endmodule

