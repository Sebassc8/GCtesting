
module cordic_DEC2_FRAC30_MOD1_DIR0 ( clk, rst, g_init, e_init, o, terminate
 );
  input [63:0] g_init;
  input [63:0] e_init;
  output [95:0] o;
  input clk, rst;
  output terminate;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N97, N98, N103, N104, N105, N106, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n508, n510, n512, n514, n516,
         n518, \add_181/carry[5] , \add_181/carry[4] , \add_181/carry[3] ,
         \add_181/carry[2] , \sub_118/carry[31] , \sub_118/carry[30] ,
         \sub_118/carry[29] , \sub_118/carry[28] , \sub_118/carry[27] ,
         \sub_118/carry[26] , \sub_118/carry[25] , \sub_118/carry[24] ,
         \sub_118/carry[23] , \sub_118/carry[22] , \sub_118/carry[21] ,
         \sub_118/carry[20] , \sub_118/carry[19] , \sub_118/carry[18] ,
         \sub_118/carry[17] , \sub_118/carry[16] , \sub_118/carry[15] ,
         \sub_118/carry[14] , \sub_118/carry[13] , \sub_118/carry[12] ,
         \sub_118/carry[11] , \sub_118/carry[10] , \sub_118/carry[9] ,
         \sub_118/carry[8] , \sub_118/carry[7] , \sub_118/carry[6] ,
         \sub_118/carry[5] , \sub_118/carry[4] , \sub_118/carry[3] ,
         \sub_118/carry[2] , \sub_115/carry[31] , \sub_115/carry[30] ,
         \sub_115/carry[29] , \sub_115/carry[28] , \sub_115/carry[27] ,
         \sub_115/carry[26] , \sub_115/carry[25] , \sub_115/carry[24] ,
         \sub_115/carry[23] , \sub_115/carry[22] , \sub_115/carry[21] ,
         \sub_115/carry[20] , \sub_115/carry[19] , \sub_115/carry[18] ,
         \sub_115/carry[17] , \sub_115/carry[16] , \sub_115/carry[15] ,
         \sub_115/carry[14] , \sub_115/carry[13] , \sub_115/carry[12] ,
         \sub_115/carry[11] , \sub_115/carry[10] , \sub_115/carry[9] ,
         \sub_115/carry[8] , \sub_115/carry[7] , \sub_115/carry[6] ,
         \sub_115/carry[5] , \sub_115/carry[4] , \sub_115/carry[3] ,
         \sub_115/carry[2] , \sub_109/carry[30] , \sub_109/carry[29] ,
         \sub_109/carry[28] , \sub_109/carry[27] , \sub_109/carry[26] ,
         \sub_109/carry[25] , \sub_109/carry[24] , \sub_109/carry[23] ,
         \sub_109/carry[22] , \sub_109/carry[21] , \sub_109/carry[20] ,
         \sub_109/carry[19] , \sub_109/carry[18] , \sub_109/carry[17] ,
         \sub_109/carry[16] , \sub_109/carry[15] , \sub_109/carry[14] ,
         \sub_109/carry[13] , \sub_109/carry[12] , \sub_109/carry[11] ,
         \sub_109/carry[10] , \sub_109/carry[9] , \sub_109/carry[8] ,
         \sub_109/carry[7] , \sub_109/carry[6] , \sub_109/carry[5] ,
         \sub_109/carry[4] , \sub_109/carry[3] , \sub_109/carry[2] , n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618;
  wire   [5:0] iter;

  DFF \iter_reg[0]  ( .D(n518), .CLK(clk), .RST(rst), .I(1'b0), .Q(iter[0]) );
  DFF \iter_reg[5]  ( .D(n516), .CLK(clk), .RST(rst), .I(1'b0), .Q(iter[5]) );
  DFF \iter_reg[1]  ( .D(n514), .CLK(clk), .RST(rst), .I(1'b0), .Q(iter[1]) );
  DFF \iter_reg[2]  ( .D(n512), .CLK(clk), .RST(rst), .I(1'b0), .Q(iter[2]) );
  DFF \iter_reg[3]  ( .D(n510), .CLK(clk), .RST(rst), .I(1'b0), .Q(iter[3]) );
  DFF \iter_reg[4]  ( .D(n508), .CLK(clk), .RST(rst), .I(1'b0), .Q(iter[4]) );
  DFF \zi_reg[28]  ( .D(n506), .CLK(clk), .RST(rst), .I(e_init[28]), .Q(o[28])
         );
  DFF \zi_reg[0]  ( .D(n505), .CLK(clk), .RST(rst), .I(e_init[0]), .Q(o[0]) );
  DFF \zi_reg[1]  ( .D(n504), .CLK(clk), .RST(rst), .I(e_init[1]), .Q(o[1]) );
  DFF \zi_reg[2]  ( .D(n503), .CLK(clk), .RST(rst), .I(e_init[2]), .Q(o[2]) );
  DFF \zi_reg[3]  ( .D(n502), .CLK(clk), .RST(rst), .I(e_init[3]), .Q(o[3]) );
  DFF \zi_reg[4]  ( .D(n501), .CLK(clk), .RST(rst), .I(e_init[4]), .Q(o[4]) );
  DFF \zi_reg[5]  ( .D(n500), .CLK(clk), .RST(rst), .I(e_init[5]), .Q(o[5]) );
  DFF \zi_reg[6]  ( .D(n499), .CLK(clk), .RST(rst), .I(e_init[6]), .Q(o[6]) );
  DFF \zi_reg[7]  ( .D(n498), .CLK(clk), .RST(rst), .I(e_init[7]), .Q(o[7]) );
  DFF \zi_reg[8]  ( .D(n497), .CLK(clk), .RST(rst), .I(e_init[8]), .Q(o[8]) );
  DFF \zi_reg[9]  ( .D(n496), .CLK(clk), .RST(rst), .I(e_init[9]), .Q(o[9]) );
  DFF \zi_reg[10]  ( .D(n495), .CLK(clk), .RST(rst), .I(e_init[10]), .Q(o[10])
         );
  DFF \zi_reg[11]  ( .D(n494), .CLK(clk), .RST(rst), .I(e_init[11]), .Q(o[11])
         );
  DFF \zi_reg[12]  ( .D(n493), .CLK(clk), .RST(rst), .I(e_init[12]), .Q(o[12])
         );
  DFF \zi_reg[13]  ( .D(n492), .CLK(clk), .RST(rst), .I(e_init[13]), .Q(o[13])
         );
  DFF \zi_reg[14]  ( .D(n491), .CLK(clk), .RST(rst), .I(e_init[14]), .Q(o[14])
         );
  DFF \zi_reg[15]  ( .D(n490), .CLK(clk), .RST(rst), .I(e_init[15]), .Q(o[15])
         );
  DFF \zi_reg[16]  ( .D(n489), .CLK(clk), .RST(rst), .I(e_init[16]), .Q(o[16])
         );
  DFF \zi_reg[17]  ( .D(n488), .CLK(clk), .RST(rst), .I(e_init[17]), .Q(o[17])
         );
  DFF \zi_reg[18]  ( .D(n487), .CLK(clk), .RST(rst), .I(e_init[18]), .Q(o[18])
         );
  DFF \zi_reg[19]  ( .D(n486), .CLK(clk), .RST(rst), .I(e_init[19]), .Q(o[19])
         );
  DFF \zi_reg[20]  ( .D(n485), .CLK(clk), .RST(rst), .I(e_init[20]), .Q(o[20])
         );
  DFF \zi_reg[21]  ( .D(n484), .CLK(clk), .RST(rst), .I(e_init[21]), .Q(o[21])
         );
  DFF \zi_reg[22]  ( .D(n483), .CLK(clk), .RST(rst), .I(e_init[22]), .Q(o[22])
         );
  DFF \zi_reg[23]  ( .D(n482), .CLK(clk), .RST(rst), .I(e_init[23]), .Q(o[23])
         );
  DFF \zi_reg[24]  ( .D(n481), .CLK(clk), .RST(rst), .I(e_init[24]), .Q(o[24])
         );
  DFF \zi_reg[25]  ( .D(n480), .CLK(clk), .RST(rst), .I(e_init[25]), .Q(o[25])
         );
  DFF \zi_reg[26]  ( .D(n479), .CLK(clk), .RST(rst), .I(e_init[26]), .Q(o[26])
         );
  DFF \zi_reg[27]  ( .D(n478), .CLK(clk), .RST(rst), .I(e_init[27]), .Q(o[27])
         );
  DFF \zi_reg[29]  ( .D(n477), .CLK(clk), .RST(rst), .I(e_init[29]), .Q(o[29])
         );
  DFF \zi_reg[30]  ( .D(n476), .CLK(clk), .RST(rst), .I(e_init[30]), .Q(o[30])
         );
  DFF \zi_reg[31]  ( .D(n475), .CLK(clk), .RST(rst), .I(e_init[31]), .Q(o[31])
         );
  DFF \yi_reg[0]  ( .D(n474), .CLK(clk), .RST(rst), .I(g_init[0]), .Q(o[32])
         );
  DFF \yi_reg[1]  ( .D(n473), .CLK(clk), .RST(rst), .I(g_init[1]), .Q(o[33])
         );
  DFF \yi_reg[2]  ( .D(n472), .CLK(clk), .RST(rst), .I(g_init[2]), .Q(o[34])
         );
  DFF \yi_reg[3]  ( .D(n471), .CLK(clk), .RST(rst), .I(g_init[3]), .Q(o[35])
         );
  DFF \yi_reg[4]  ( .D(n470), .CLK(clk), .RST(rst), .I(g_init[4]), .Q(o[36])
         );
  DFF \yi_reg[5]  ( .D(n469), .CLK(clk), .RST(rst), .I(g_init[5]), .Q(o[37])
         );
  DFF \yi_reg[6]  ( .D(n468), .CLK(clk), .RST(rst), .I(g_init[6]), .Q(o[38])
         );
  DFF \yi_reg[7]  ( .D(n467), .CLK(clk), .RST(rst), .I(g_init[7]), .Q(o[39])
         );
  DFF \yi_reg[8]  ( .D(n466), .CLK(clk), .RST(rst), .I(g_init[8]), .Q(o[40])
         );
  DFF \yi_reg[9]  ( .D(n465), .CLK(clk), .RST(rst), .I(g_init[9]), .Q(o[41])
         );
  DFF \yi_reg[10]  ( .D(n464), .CLK(clk), .RST(rst), .I(g_init[10]), .Q(o[42])
         );
  DFF \yi_reg[11]  ( .D(n463), .CLK(clk), .RST(rst), .I(g_init[11]), .Q(o[43])
         );
  DFF \yi_reg[12]  ( .D(n462), .CLK(clk), .RST(rst), .I(g_init[12]), .Q(o[44])
         );
  DFF \yi_reg[13]  ( .D(n461), .CLK(clk), .RST(rst), .I(g_init[13]), .Q(o[45])
         );
  DFF \yi_reg[14]  ( .D(n460), .CLK(clk), .RST(rst), .I(g_init[14]), .Q(o[46])
         );
  DFF \yi_reg[15]  ( .D(n459), .CLK(clk), .RST(rst), .I(g_init[15]), .Q(o[47])
         );
  DFF \yi_reg[16]  ( .D(n458), .CLK(clk), .RST(rst), .I(g_init[16]), .Q(o[48])
         );
  DFF \yi_reg[17]  ( .D(n457), .CLK(clk), .RST(rst), .I(g_init[17]), .Q(o[49])
         );
  DFF \yi_reg[18]  ( .D(n456), .CLK(clk), .RST(rst), .I(g_init[18]), .Q(o[50])
         );
  DFF \yi_reg[19]  ( .D(n455), .CLK(clk), .RST(rst), .I(g_init[19]), .Q(o[51])
         );
  DFF \yi_reg[20]  ( .D(n454), .CLK(clk), .RST(rst), .I(g_init[20]), .Q(o[52])
         );
  DFF \yi_reg[21]  ( .D(n453), .CLK(clk), .RST(rst), .I(g_init[21]), .Q(o[53])
         );
  DFF \yi_reg[22]  ( .D(n452), .CLK(clk), .RST(rst), .I(g_init[22]), .Q(o[54])
         );
  DFF \yi_reg[23]  ( .D(n451), .CLK(clk), .RST(rst), .I(g_init[23]), .Q(o[55])
         );
  DFF \yi_reg[24]  ( .D(n450), .CLK(clk), .RST(rst), .I(g_init[24]), .Q(o[56])
         );
  DFF \yi_reg[25]  ( .D(n449), .CLK(clk), .RST(rst), .I(g_init[25]), .Q(o[57])
         );
  DFF \yi_reg[26]  ( .D(n448), .CLK(clk), .RST(rst), .I(g_init[26]), .Q(o[58])
         );
  DFF \yi_reg[27]  ( .D(n447), .CLK(clk), .RST(rst), .I(g_init[27]), .Q(o[59])
         );
  DFF \yi_reg[28]  ( .D(n446), .CLK(clk), .RST(rst), .I(g_init[28]), .Q(o[60])
         );
  DFF \yi_reg[29]  ( .D(n445), .CLK(clk), .RST(rst), .I(g_init[29]), .Q(o[61])
         );
  DFF \yi_reg[30]  ( .D(n444), .CLK(clk), .RST(rst), .I(g_init[30]), .Q(o[62])
         );
  DFF \yi_reg[31]  ( .D(n443), .CLK(clk), .RST(rst), .I(g_init[31]), .Q(o[63])
         );
  DFF \xi_reg[0]  ( .D(n442), .CLK(clk), .RST(rst), .I(g_init[32]), .Q(o[64])
         );
  DFF \xi_reg[1]  ( .D(n441), .CLK(clk), .RST(rst), .I(g_init[33]), .Q(o[65])
         );
  DFF \xi_reg[2]  ( .D(n440), .CLK(clk), .RST(rst), .I(g_init[34]), .Q(o[66])
         );
  DFF \xi_reg[3]  ( .D(n439), .CLK(clk), .RST(rst), .I(g_init[35]), .Q(o[67])
         );
  DFF \xi_reg[4]  ( .D(n438), .CLK(clk), .RST(rst), .I(g_init[36]), .Q(o[68])
         );
  DFF \xi_reg[5]  ( .D(n437), .CLK(clk), .RST(rst), .I(g_init[37]), .Q(o[69])
         );
  DFF \xi_reg[6]  ( .D(n436), .CLK(clk), .RST(rst), .I(g_init[38]), .Q(o[70])
         );
  DFF \xi_reg[7]  ( .D(n435), .CLK(clk), .RST(rst), .I(g_init[39]), .Q(o[71])
         );
  DFF \xi_reg[8]  ( .D(n434), .CLK(clk), .RST(rst), .I(g_init[40]), .Q(o[72])
         );
  DFF \xi_reg[9]  ( .D(n433), .CLK(clk), .RST(rst), .I(g_init[41]), .Q(o[73])
         );
  DFF \xi_reg[10]  ( .D(n432), .CLK(clk), .RST(rst), .I(g_init[42]), .Q(o[74])
         );
  DFF \xi_reg[11]  ( .D(n431), .CLK(clk), .RST(rst), .I(g_init[43]), .Q(o[75])
         );
  DFF \xi_reg[12]  ( .D(n430), .CLK(clk), .RST(rst), .I(g_init[44]), .Q(o[76])
         );
  DFF \xi_reg[13]  ( .D(n429), .CLK(clk), .RST(rst), .I(g_init[45]), .Q(o[77])
         );
  DFF \xi_reg[14]  ( .D(n428), .CLK(clk), .RST(rst), .I(g_init[46]), .Q(o[78])
         );
  DFF \xi_reg[15]  ( .D(n427), .CLK(clk), .RST(rst), .I(g_init[47]), .Q(o[79])
         );
  DFF \xi_reg[16]  ( .D(n426), .CLK(clk), .RST(rst), .I(g_init[48]), .Q(o[80])
         );
  DFF \xi_reg[17]  ( .D(n425), .CLK(clk), .RST(rst), .I(g_init[49]), .Q(o[81])
         );
  DFF \xi_reg[18]  ( .D(n424), .CLK(clk), .RST(rst), .I(g_init[50]), .Q(o[82])
         );
  DFF \xi_reg[19]  ( .D(n423), .CLK(clk), .RST(rst), .I(g_init[51]), .Q(o[83])
         );
  DFF \xi_reg[20]  ( .D(n422), .CLK(clk), .RST(rst), .I(g_init[52]), .Q(o[84])
         );
  DFF \xi_reg[21]  ( .D(n421), .CLK(clk), .RST(rst), .I(g_init[53]), .Q(o[85])
         );
  DFF \xi_reg[22]  ( .D(n420), .CLK(clk), .RST(rst), .I(g_init[54]), .Q(o[86])
         );
  DFF \xi_reg[23]  ( .D(n419), .CLK(clk), .RST(rst), .I(g_init[55]), .Q(o[87])
         );
  DFF \xi_reg[24]  ( .D(n418), .CLK(clk), .RST(rst), .I(g_init[56]), .Q(o[88])
         );
  DFF \xi_reg[25]  ( .D(n417), .CLK(clk), .RST(rst), .I(g_init[57]), .Q(o[89])
         );
  DFF \xi_reg[26]  ( .D(n416), .CLK(clk), .RST(rst), .I(g_init[58]), .Q(o[90])
         );
  DFF \xi_reg[27]  ( .D(n415), .CLK(clk), .RST(rst), .I(g_init[59]), .Q(o[91])
         );
  DFF \xi_reg[28]  ( .D(n414), .CLK(clk), .RST(rst), .I(g_init[60]), .Q(o[92])
         );
  DFF \xi_reg[29]  ( .D(n413), .CLK(clk), .RST(rst), .I(g_init[61]), .Q(o[93])
         );
  DFF \xi_reg[30]  ( .D(n412), .CLK(clk), .RST(rst), .I(g_init[62]), .Q(o[94])
         );
  DFF \xi_reg[31]  ( .D(n411), .CLK(clk), .RST(rst), .I(g_init[63]), .Q(o[95])
         );
  HADDER \add_181/U1_1_1  ( .IN0(iter[1]), .IN1(iter[0]), .COUT(
        \add_181/carry[2] ), .SUM(N103) );
  HADDER \add_181/U1_1_2  ( .IN0(iter[2]), .IN1(\add_181/carry[2] ), .COUT(
        \add_181/carry[3] ), .SUM(N104) );
  HADDER \add_181/U1_1_3  ( .IN0(iter[3]), .IN1(\add_181/carry[3] ), .COUT(
        \add_181/carry[4] ), .SUM(N105) );
  HADDER \add_181/U1_1_4  ( .IN0(iter[4]), .IN1(\add_181/carry[4] ), .COUT(
        \add_181/carry[5] ), .SUM(N106) );
  MUX U614 ( .IN0(n708), .IN1(o[26]), .SEL(n677), .F(n701) );
  MUX U615 ( .IN0(n793), .IN1(o[13]), .SEL(n651), .F(n787) );
  MUX U616 ( .IN0(n1318), .IN1(o[92]), .SEL(n1294), .F(n1315) );
  MUX U617 ( .IN0(n1330), .IN1(o[88]), .SEL(n1286), .F(n1327) );
  MUX U618 ( .IN0(n1342), .IN1(o[84]), .SEL(n1278), .F(n1339) );
  MUX U619 ( .IN0(n1354), .IN1(o[80]), .SEL(n1270), .F(n1351) );
  MUX U620 ( .IN0(n1378), .IN1(o[76]), .SEL(n1262), .F(n1371) );
  MUX U621 ( .IN0(n1406), .IN1(o[72]), .SEL(n1251), .F(n1399) );
  MUX U622 ( .IN0(n1451), .IN1(o[68]), .SEL(n1239), .F(n1439) );
  MUX U623 ( .IN0(n1006), .IN1(o[60]), .SEL(n985), .F(n1003) );
  MUX U624 ( .IN0(n1018), .IN1(o[56]), .SEL(n977), .F(n1015) );
  MUX U625 ( .IN0(n1030), .IN1(o[52]), .SEL(n969), .F(n1027) );
  MUX U626 ( .IN0(n1042), .IN1(o[48]), .SEL(n961), .F(n1039) );
  MUX U627 ( .IN0(n1066), .IN1(o[44]), .SEL(n953), .F(n1059) );
  MUX U628 ( .IN0(n1094), .IN1(o[40]), .SEL(n939), .F(n1087) );
  MUX U629 ( .IN0(n1139), .IN1(o[36]), .SEL(n923), .F(n1127) );
  MUX U630 ( .IN0(n712), .IN1(o[25]), .SEL(n675), .F(n708) );
  MUX U631 ( .IN0(n737), .IN1(o[21]), .SEL(n667), .F(n730) );
  MUX U632 ( .IN0(n769), .IN1(o[17]), .SEL(n659), .F(n764) );
  MUX U633 ( .IN0(n802), .IN1(o[12]), .SEL(n649), .F(n793) );
  MUX U634 ( .IN0(n830), .IN1(o[8]), .SEL(n641), .F(n824) );
  MUX U635 ( .IN0(n857), .IN1(o[4]), .SEL(n633), .F(n852) );
  MUX U636 ( .IN0(n1321), .IN1(o[91]), .SEL(n1292), .F(n1318) );
  MUX U637 ( .IN0(n1333), .IN1(o[87]), .SEL(n1284), .F(n1330) );
  MUX U638 ( .IN0(n1345), .IN1(o[83]), .SEL(n1276), .F(n1342) );
  MUX U639 ( .IN0(n1357), .IN1(o[79]), .SEL(n1268), .F(n1354) );
  MUX U640 ( .IN0(n1385), .IN1(o[75]), .SEL(n1260), .F(n1378) );
  MUX U641 ( .IN0(n1413), .IN1(o[71]), .SEL(n1248), .F(n1406) );
  MUX U642 ( .IN0(n1465), .IN1(o[67]), .SEL(n1236), .F(n1451) );
  MUX U643 ( .IN0(n1009), .IN1(o[59]), .SEL(n983), .F(n1006) );
  MUX U644 ( .IN0(n1021), .IN1(o[55]), .SEL(n975), .F(n1018) );
  MUX U645 ( .IN0(n1033), .IN1(o[51]), .SEL(n967), .F(n1030) );
  MUX U646 ( .IN0(n1045), .IN1(o[47]), .SEL(n959), .F(n1042) );
  MUX U647 ( .IN0(n1073), .IN1(o[43]), .SEL(n951), .F(n1066) );
  MUX U648 ( .IN0(n1101), .IN1(o[39]), .SEL(n935), .F(n1094) );
  MUX U649 ( .IN0(n1153), .IN1(o[35]), .SEL(n919), .F(n1139) );
  MUX U650 ( .IN0(n694), .IN1(o[29]), .SEL(n681), .F(n520) );
  IV U651 ( .A(n520), .Z(n693) );
  MUX U652 ( .IN0(n715), .IN1(o[24]), .SEL(n673), .F(n712) );
  MUX U653 ( .IN0(n744), .IN1(o[20]), .SEL(n665), .F(n737) );
  MUX U654 ( .IN0(n773), .IN1(o[16]), .SEL(n657), .F(n769) );
  MUX U655 ( .IN0(n810), .IN1(o[11]), .SEL(n647), .F(n802) );
  MUX U656 ( .IN0(n837), .IN1(o[7]), .SEL(n639), .F(n830) );
  MUX U657 ( .IN0(n868), .IN1(o[3]), .SEL(n631), .F(n857) );
  ANDN U658 ( .A(n777), .B(n734), .Z(n766) );
  MUX U659 ( .IN0(n1324), .IN1(o[90]), .SEL(n1290), .F(n1321) );
  MUX U660 ( .IN0(n1336), .IN1(o[86]), .SEL(n1282), .F(n1333) );
  MUX U661 ( .IN0(n1348), .IN1(o[82]), .SEL(n1274), .F(n1345) );
  MUX U662 ( .IN0(n1364), .IN1(o[78]), .SEL(n1266), .F(n1357) );
  MUX U663 ( .IN0(n1392), .IN1(o[74]), .SEL(n1257), .F(n1385) );
  MUX U664 ( .IN0(n1425), .IN1(o[70]), .SEL(n1245), .F(n1413) );
  MUX U665 ( .IN0(n1487), .IN1(o[66]), .SEL(n1233), .F(n1465) );
  MUX U666 ( .IN0(n1012), .IN1(o[58]), .SEL(n981), .F(n1009) );
  MUX U667 ( .IN0(n1024), .IN1(o[54]), .SEL(n973), .F(n1021) );
  MUX U668 ( .IN0(n1036), .IN1(o[50]), .SEL(n965), .F(n1033) );
  MUX U669 ( .IN0(n1052), .IN1(o[46]), .SEL(n957), .F(n1045) );
  MUX U670 ( .IN0(n1080), .IN1(o[42]), .SEL(n947), .F(n1073) );
  MUX U671 ( .IN0(n1113), .IN1(o[38]), .SEL(n931), .F(n1101) );
  MUX U672 ( .IN0(n1175), .IN1(o[34]), .SEL(n915), .F(n1153) );
  MUX U673 ( .IN0(n697), .IN1(o[28]), .SEL(n624), .F(n694) );
  MUX U674 ( .IN0(n719), .IN1(o[23]), .SEL(n671), .F(n715) );
  MUX U675 ( .IN0(n750), .IN1(o[19]), .SEL(n663), .F(n744) );
  MUX U676 ( .IN0(n783), .IN1(o[15]), .SEL(n655), .F(n773) );
  MUX U677 ( .IN0(n819), .IN1(o[10]), .SEL(n645), .F(n810) );
  MUX U678 ( .IN0(n847), .IN1(o[6]), .SEL(n637), .F(n837) );
  MUX U679 ( .IN0(n876), .IN1(o[2]), .SEL(n629), .F(n868) );
  XNOR U680 ( .A(n552), .B(\sub_115/carry[31] ), .Z(N66) );
  XNOR U681 ( .A(n583), .B(\sub_118/carry[31] ), .Z(N98) );
  MUX U682 ( .IN0(n1327), .IN1(o[89]), .SEL(n1288), .F(n1324) );
  MUX U683 ( .IN0(n1339), .IN1(o[85]), .SEL(n1280), .F(n1336) );
  MUX U684 ( .IN0(n1351), .IN1(o[81]), .SEL(n1272), .F(n1348) );
  MUX U685 ( .IN0(n1371), .IN1(o[77]), .SEL(n1264), .F(n1364) );
  MUX U686 ( .IN0(n1399), .IN1(o[73]), .SEL(n1254), .F(n1392) );
  MUX U687 ( .IN0(n1439), .IN1(o[69]), .SEL(n1242), .F(n1425) );
  MUX U688 ( .IN0(o[65]), .IN1(n521), .SEL(n1230), .F(n1487) );
  IV U689 ( .A(n1512), .Z(n521) );
  MUX U690 ( .IN0(n1015), .IN1(o[57]), .SEL(n979), .F(n1012) );
  MUX U691 ( .IN0(n1027), .IN1(o[53]), .SEL(n971), .F(n1024) );
  MUX U692 ( .IN0(n1039), .IN1(o[49]), .SEL(n963), .F(n1036) );
  MUX U693 ( .IN0(n1059), .IN1(o[45]), .SEL(n955), .F(n1052) );
  MUX U694 ( .IN0(n1087), .IN1(o[41]), .SEL(n943), .F(n1080) );
  MUX U695 ( .IN0(n1127), .IN1(o[37]), .SEL(n927), .F(n1113) );
  MUX U696 ( .IN0(o[33]), .IN1(n522), .SEL(n911), .F(n1175) );
  IV U697 ( .A(n1200), .Z(n522) );
  MUX U698 ( .IN0(n730), .IN1(o[22]), .SEL(n669), .F(n719) );
  MUX U699 ( .IN0(n764), .IN1(o[18]), .SEL(n661), .F(n750) );
  MUX U700 ( .IN0(n787), .IN1(o[14]), .SEL(n653), .F(n783) );
  NANDN U701 ( .B(n736), .A(n801), .Z(n800) );
  MUX U702 ( .IN0(n824), .IN1(o[9]), .SEL(n643), .F(n819) );
  MUX U703 ( .IN0(n852), .IN1(o[5]), .SEL(n635), .F(n847) );
  MUX U704 ( .IN0(n890), .IN1(o[1]), .SEL(n627), .F(n876) );
  MUX U705 ( .IN0(n701), .IN1(o[27]), .SEL(n679), .F(n697) );
  MUX U706 ( .IN0(n1315), .IN1(o[93]), .SEL(n1296), .F(n1308) );
  MUX U707 ( .IN0(n1003), .IN1(o[61]), .SEL(n987), .F(n995) );
  AND U708 ( .A(n1586), .B(n1558), .Z(\sub_118/carry[2] ) );
  XOR U709 ( .A(n1586), .B(n1558), .Z(N68) );
  AND U710 ( .A(n1569), .B(\sub_118/carry[2] ), .Z(\sub_118/carry[3] ) );
  XOR U711 ( .A(n1569), .B(\sub_118/carry[2] ), .Z(N69) );
  AND U712 ( .A(n1577), .B(\sub_118/carry[3] ), .Z(\sub_118/carry[4] ) );
  XOR U713 ( .A(n1577), .B(\sub_118/carry[3] ), .Z(N70) );
  AND U714 ( .A(n1565), .B(\sub_118/carry[4] ), .Z(\sub_118/carry[5] ) );
  XOR U715 ( .A(n1565), .B(\sub_118/carry[4] ), .Z(N71) );
  AND U716 ( .A(n1584), .B(\sub_118/carry[5] ), .Z(\sub_118/carry[6] ) );
  XOR U717 ( .A(n1584), .B(\sub_118/carry[5] ), .Z(N72) );
  AND U718 ( .A(n1573), .B(\sub_118/carry[6] ), .Z(\sub_118/carry[7] ) );
  XOR U719 ( .A(n1573), .B(\sub_118/carry[6] ), .Z(N73) );
  AND U720 ( .A(n1580), .B(\sub_118/carry[7] ), .Z(\sub_118/carry[8] ) );
  XOR U721 ( .A(n1580), .B(\sub_118/carry[7] ), .Z(N74) );
  AND U722 ( .A(n1561), .B(\sub_118/carry[8] ), .Z(\sub_118/carry[9] ) );
  XOR U723 ( .A(n1561), .B(\sub_118/carry[8] ), .Z(N75) );
  AND U724 ( .A(n1588), .B(\sub_118/carry[9] ), .Z(\sub_118/carry[10] ) );
  XOR U725 ( .A(n1588), .B(\sub_118/carry[9] ), .Z(N76) );
  AND U726 ( .A(n1566), .B(\sub_118/carry[10] ), .Z(\sub_118/carry[11] ) );
  XOR U727 ( .A(n1566), .B(\sub_118/carry[10] ), .Z(N77) );
  AND U728 ( .A(n1574), .B(\sub_118/carry[11] ), .Z(\sub_118/carry[12] ) );
  XOR U729 ( .A(n1574), .B(\sub_118/carry[11] ), .Z(N78) );
  AND U730 ( .A(n1562), .B(\sub_118/carry[12] ), .Z(\sub_118/carry[13] ) );
  XOR U731 ( .A(n1562), .B(\sub_118/carry[12] ), .Z(N79) );
  AND U732 ( .A(n1581), .B(\sub_118/carry[13] ), .Z(\sub_118/carry[14] ) );
  XOR U733 ( .A(n1581), .B(\sub_118/carry[13] ), .Z(N80) );
  AND U734 ( .A(n1570), .B(\sub_118/carry[14] ), .Z(\sub_118/carry[15] ) );
  XOR U735 ( .A(n1570), .B(\sub_118/carry[14] ), .Z(N81) );
  AND U736 ( .A(n1578), .B(\sub_118/carry[15] ), .Z(\sub_118/carry[16] ) );
  XOR U737 ( .A(n1578), .B(\sub_118/carry[15] ), .Z(N82) );
  AND U738 ( .A(n1559), .B(\sub_118/carry[16] ), .Z(\sub_118/carry[17] ) );
  XOR U739 ( .A(n1559), .B(\sub_118/carry[16] ), .Z(N83) );
  AND U740 ( .A(n1585), .B(\sub_118/carry[17] ), .Z(\sub_118/carry[18] ) );
  XOR U741 ( .A(n1585), .B(\sub_118/carry[17] ), .Z(N84) );
  AND U742 ( .A(n1568), .B(\sub_118/carry[18] ), .Z(\sub_118/carry[19] ) );
  XOR U743 ( .A(n1568), .B(\sub_118/carry[18] ), .Z(N85) );
  AND U744 ( .A(n1576), .B(\sub_118/carry[19] ), .Z(\sub_118/carry[20] ) );
  XOR U745 ( .A(n1576), .B(\sub_118/carry[19] ), .Z(N86) );
  AND U746 ( .A(n1564), .B(\sub_118/carry[20] ), .Z(\sub_118/carry[21] ) );
  XOR U747 ( .A(n1564), .B(\sub_118/carry[20] ), .Z(N87) );
  AND U748 ( .A(n1583), .B(\sub_118/carry[21] ), .Z(\sub_118/carry[22] ) );
  XOR U749 ( .A(n1583), .B(\sub_118/carry[21] ), .Z(N88) );
  AND U750 ( .A(n1572), .B(\sub_118/carry[22] ), .Z(\sub_118/carry[23] ) );
  XOR U751 ( .A(n1572), .B(\sub_118/carry[22] ), .Z(N89) );
  AND U752 ( .A(n1579), .B(\sub_118/carry[23] ), .Z(\sub_118/carry[24] ) );
  XOR U753 ( .A(n1579), .B(\sub_118/carry[23] ), .Z(N90) );
  AND U754 ( .A(n1560), .B(\sub_118/carry[24] ), .Z(\sub_118/carry[25] ) );
  XOR U755 ( .A(n1560), .B(\sub_118/carry[24] ), .Z(N91) );
  AND U756 ( .A(n1587), .B(\sub_118/carry[25] ), .Z(\sub_118/carry[26] ) );
  XOR U757 ( .A(n1587), .B(\sub_118/carry[25] ), .Z(N92) );
  AND U758 ( .A(n1567), .B(\sub_118/carry[26] ), .Z(\sub_118/carry[27] ) );
  XOR U759 ( .A(n1567), .B(\sub_118/carry[26] ), .Z(N93) );
  AND U760 ( .A(n1575), .B(\sub_118/carry[27] ), .Z(\sub_118/carry[28] ) );
  XOR U761 ( .A(n1575), .B(\sub_118/carry[27] ), .Z(N94) );
  AND U762 ( .A(n1563), .B(\sub_118/carry[28] ), .Z(\sub_118/carry[29] ) );
  XOR U763 ( .A(n1563), .B(\sub_118/carry[28] ), .Z(N95) );
  AND U764 ( .A(n1582), .B(\sub_118/carry[29] ), .Z(\sub_118/carry[30] ) );
  XOR U765 ( .A(n1582), .B(\sub_118/carry[29] ), .Z(N96) );
  AND U766 ( .A(n1571), .B(\sub_118/carry[30] ), .Z(\sub_118/carry[31] ) );
  XOR U767 ( .A(n1571), .B(\sub_118/carry[30] ), .Z(N97) );
  AND U768 ( .A(n1555), .B(n1527), .Z(\sub_115/carry[2] ) );
  XOR U769 ( .A(n1555), .B(n1527), .Z(N36) );
  AND U770 ( .A(n1538), .B(\sub_115/carry[2] ), .Z(\sub_115/carry[3] ) );
  XOR U771 ( .A(n1538), .B(\sub_115/carry[2] ), .Z(N37) );
  AND U772 ( .A(n1546), .B(\sub_115/carry[3] ), .Z(\sub_115/carry[4] ) );
  XOR U773 ( .A(n1546), .B(\sub_115/carry[3] ), .Z(N38) );
  AND U774 ( .A(n1534), .B(\sub_115/carry[4] ), .Z(\sub_115/carry[5] ) );
  XOR U775 ( .A(n1534), .B(\sub_115/carry[4] ), .Z(N39) );
  AND U776 ( .A(n1553), .B(\sub_115/carry[5] ), .Z(\sub_115/carry[6] ) );
  XOR U777 ( .A(n1553), .B(\sub_115/carry[5] ), .Z(N40) );
  AND U778 ( .A(n1542), .B(\sub_115/carry[6] ), .Z(\sub_115/carry[7] ) );
  XOR U779 ( .A(n1542), .B(\sub_115/carry[6] ), .Z(N41) );
  AND U780 ( .A(n1549), .B(\sub_115/carry[7] ), .Z(\sub_115/carry[8] ) );
  XOR U781 ( .A(n1549), .B(\sub_115/carry[7] ), .Z(N42) );
  AND U782 ( .A(n1530), .B(\sub_115/carry[8] ), .Z(\sub_115/carry[9] ) );
  XOR U783 ( .A(n1530), .B(\sub_115/carry[8] ), .Z(N43) );
  AND U784 ( .A(n1557), .B(\sub_115/carry[9] ), .Z(\sub_115/carry[10] ) );
  XOR U785 ( .A(n1557), .B(\sub_115/carry[9] ), .Z(N44) );
  AND U786 ( .A(n1535), .B(\sub_115/carry[10] ), .Z(\sub_115/carry[11] ) );
  XOR U787 ( .A(n1535), .B(\sub_115/carry[10] ), .Z(N45) );
  AND U788 ( .A(n1543), .B(\sub_115/carry[11] ), .Z(\sub_115/carry[12] ) );
  XOR U789 ( .A(n1543), .B(\sub_115/carry[11] ), .Z(N46) );
  AND U790 ( .A(n1531), .B(\sub_115/carry[12] ), .Z(\sub_115/carry[13] ) );
  XOR U791 ( .A(n1531), .B(\sub_115/carry[12] ), .Z(N47) );
  AND U792 ( .A(n1550), .B(\sub_115/carry[13] ), .Z(\sub_115/carry[14] ) );
  XOR U793 ( .A(n1550), .B(\sub_115/carry[13] ), .Z(N48) );
  AND U794 ( .A(n1539), .B(\sub_115/carry[14] ), .Z(\sub_115/carry[15] ) );
  XOR U795 ( .A(n1539), .B(\sub_115/carry[14] ), .Z(N49) );
  AND U796 ( .A(n1547), .B(\sub_115/carry[15] ), .Z(\sub_115/carry[16] ) );
  XOR U797 ( .A(n1547), .B(\sub_115/carry[15] ), .Z(N50) );
  AND U798 ( .A(n1528), .B(\sub_115/carry[16] ), .Z(\sub_115/carry[17] ) );
  XOR U799 ( .A(n1528), .B(\sub_115/carry[16] ), .Z(N51) );
  AND U800 ( .A(n1554), .B(\sub_115/carry[17] ), .Z(\sub_115/carry[18] ) );
  XOR U801 ( .A(n1554), .B(\sub_115/carry[17] ), .Z(N52) );
  AND U802 ( .A(n1537), .B(\sub_115/carry[18] ), .Z(\sub_115/carry[19] ) );
  XOR U803 ( .A(n1537), .B(\sub_115/carry[18] ), .Z(N53) );
  AND U804 ( .A(n1545), .B(\sub_115/carry[19] ), .Z(\sub_115/carry[20] ) );
  XOR U805 ( .A(n1545), .B(\sub_115/carry[19] ), .Z(N54) );
  AND U806 ( .A(n1533), .B(\sub_115/carry[20] ), .Z(\sub_115/carry[21] ) );
  XOR U807 ( .A(n1533), .B(\sub_115/carry[20] ), .Z(N55) );
  AND U808 ( .A(n1552), .B(\sub_115/carry[21] ), .Z(\sub_115/carry[22] ) );
  XOR U809 ( .A(n1552), .B(\sub_115/carry[21] ), .Z(N56) );
  AND U810 ( .A(n1541), .B(\sub_115/carry[22] ), .Z(\sub_115/carry[23] ) );
  XOR U811 ( .A(n1541), .B(\sub_115/carry[22] ), .Z(N57) );
  AND U812 ( .A(n1548), .B(\sub_115/carry[23] ), .Z(\sub_115/carry[24] ) );
  XOR U813 ( .A(n1548), .B(\sub_115/carry[23] ), .Z(N58) );
  AND U814 ( .A(n1529), .B(\sub_115/carry[24] ), .Z(\sub_115/carry[25] ) );
  XOR U815 ( .A(n1529), .B(\sub_115/carry[24] ), .Z(N59) );
  AND U816 ( .A(n1556), .B(\sub_115/carry[25] ), .Z(\sub_115/carry[26] ) );
  XOR U817 ( .A(n1556), .B(\sub_115/carry[25] ), .Z(N60) );
  AND U818 ( .A(n1536), .B(\sub_115/carry[26] ), .Z(\sub_115/carry[27] ) );
  XOR U819 ( .A(n1536), .B(\sub_115/carry[26] ), .Z(N61) );
  AND U820 ( .A(n1544), .B(\sub_115/carry[27] ), .Z(\sub_115/carry[28] ) );
  XOR U821 ( .A(n1544), .B(\sub_115/carry[27] ), .Z(N62) );
  AND U822 ( .A(n1532), .B(\sub_115/carry[28] ), .Z(\sub_115/carry[29] ) );
  XOR U823 ( .A(n1532), .B(\sub_115/carry[28] ), .Z(N63) );
  AND U824 ( .A(n1551), .B(\sub_115/carry[29] ), .Z(\sub_115/carry[30] ) );
  XOR U825 ( .A(n1551), .B(\sub_115/carry[29] ), .Z(N64) );
  AND U826 ( .A(n1540), .B(\sub_115/carry[30] ), .Z(\sub_115/carry[31] ) );
  XOR U827 ( .A(n1540), .B(\sub_115/carry[30] ), .Z(N65) );
  AND U828 ( .A(n1591), .B(n1600), .Z(\sub_109/carry[2] ) );
  XOR U829 ( .A(n1591), .B(n1600), .Z(N4) );
  AND U830 ( .A(n1595), .B(\sub_109/carry[2] ), .Z(\sub_109/carry[3] ) );
  XOR U831 ( .A(n1595), .B(\sub_109/carry[2] ), .Z(N5) );
  AND U832 ( .A(n1589), .B(\sub_109/carry[3] ), .Z(\sub_109/carry[4] ) );
  XOR U833 ( .A(n1589), .B(\sub_109/carry[3] ), .Z(N6) );
  AND U834 ( .A(n1604), .B(\sub_109/carry[4] ), .Z(\sub_109/carry[5] ) );
  XOR U835 ( .A(n1604), .B(\sub_109/carry[4] ), .Z(N7) );
  AND U836 ( .A(n1611), .B(\sub_109/carry[5] ), .Z(\sub_109/carry[6] ) );
  XOR U837 ( .A(n1611), .B(\sub_109/carry[5] ), .Z(N8) );
  AND U838 ( .A(n1603), .B(\sub_109/carry[6] ), .Z(\sub_109/carry[7] ) );
  XOR U839 ( .A(n1603), .B(\sub_109/carry[6] ), .Z(N9) );
  AND U840 ( .A(n1590), .B(\sub_109/carry[7] ), .Z(\sub_109/carry[8] ) );
  XOR U841 ( .A(n1590), .B(\sub_109/carry[7] ), .Z(N10) );
  AND U842 ( .A(n1602), .B(\sub_109/carry[8] ), .Z(\sub_109/carry[9] ) );
  XOR U843 ( .A(n1602), .B(\sub_109/carry[8] ), .Z(N11) );
  AND U844 ( .A(n1610), .B(\sub_109/carry[9] ), .Z(\sub_109/carry[10] ) );
  XOR U845 ( .A(n1610), .B(\sub_109/carry[9] ), .Z(N12) );
  AND U846 ( .A(n1609), .B(\sub_109/carry[10] ), .Z(\sub_109/carry[11] ) );
  XOR U847 ( .A(n1609), .B(\sub_109/carry[10] ), .Z(N13) );
  AND U848 ( .A(n1592), .B(\sub_109/carry[11] ), .Z(\sub_109/carry[12] ) );
  XOR U849 ( .A(n1592), .B(\sub_109/carry[11] ), .Z(N14) );
  AND U850 ( .A(n1601), .B(\sub_109/carry[12] ), .Z(\sub_109/carry[13] ) );
  XOR U851 ( .A(n1601), .B(\sub_109/carry[12] ), .Z(N15) );
  AND U852 ( .A(n1599), .B(\sub_109/carry[13] ), .Z(\sub_109/carry[14] ) );
  XOR U853 ( .A(n1599), .B(\sub_109/carry[13] ), .Z(N16) );
  AND U854 ( .A(n1608), .B(\sub_109/carry[14] ), .Z(\sub_109/carry[15] ) );
  XOR U855 ( .A(n1608), .B(\sub_109/carry[14] ), .Z(N17) );
  AND U856 ( .A(n1617), .B(\sub_109/carry[15] ), .Z(\sub_109/carry[16] ) );
  XOR U857 ( .A(n1617), .B(\sub_109/carry[15] ), .Z(N18) );
  AND U858 ( .A(n1616), .B(\sub_109/carry[16] ), .Z(\sub_109/carry[17] ) );
  XOR U859 ( .A(n1616), .B(\sub_109/carry[16] ), .Z(N19) );
  AND U860 ( .A(n1607), .B(\sub_109/carry[17] ), .Z(\sub_109/carry[18] ) );
  XOR U861 ( .A(n1607), .B(\sub_109/carry[17] ), .Z(N20) );
  AND U862 ( .A(n1615), .B(\sub_109/carry[18] ), .Z(\sub_109/carry[19] ) );
  XOR U863 ( .A(n1615), .B(\sub_109/carry[18] ), .Z(N21) );
  AND U864 ( .A(n1594), .B(\sub_109/carry[19] ), .Z(\sub_109/carry[20] ) );
  XOR U865 ( .A(n1594), .B(\sub_109/carry[19] ), .Z(N22) );
  AND U866 ( .A(n1612), .B(\sub_109/carry[20] ), .Z(\sub_109/carry[21] ) );
  XOR U867 ( .A(n1612), .B(\sub_109/carry[20] ), .Z(N23) );
  AND U868 ( .A(n1593), .B(\sub_109/carry[21] ), .Z(\sub_109/carry[22] ) );
  XOR U869 ( .A(n1593), .B(\sub_109/carry[21] ), .Z(N24) );
  AND U870 ( .A(n1598), .B(\sub_109/carry[22] ), .Z(\sub_109/carry[23] ) );
  XOR U871 ( .A(n1598), .B(\sub_109/carry[22] ), .Z(N25) );
  AND U872 ( .A(n1606), .B(\sub_109/carry[23] ), .Z(\sub_109/carry[24] ) );
  XOR U873 ( .A(n1606), .B(\sub_109/carry[23] ), .Z(N26) );
  AND U874 ( .A(n1614), .B(\sub_109/carry[24] ), .Z(\sub_109/carry[25] ) );
  XOR U875 ( .A(n1614), .B(\sub_109/carry[24] ), .Z(N27) );
  AND U876 ( .A(n1597), .B(\sub_109/carry[25] ), .Z(\sub_109/carry[26] ) );
  XOR U877 ( .A(n1597), .B(\sub_109/carry[25] ), .Z(N28) );
  AND U878 ( .A(n1613), .B(\sub_109/carry[26] ), .Z(\sub_109/carry[27] ) );
  XOR U879 ( .A(n1613), .B(\sub_109/carry[26] ), .Z(N29) );
  AND U880 ( .A(n1596), .B(\sub_109/carry[27] ), .Z(\sub_109/carry[28] ) );
  XOR U881 ( .A(n1596), .B(\sub_109/carry[27] ), .Z(N30) );
  AND U882 ( .A(n1618), .B(\sub_109/carry[28] ), .Z(\sub_109/carry[29] ) );
  XOR U883 ( .A(n1618), .B(\sub_109/carry[28] ), .Z(N31) );
  AND U884 ( .A(n1605), .B(\sub_109/carry[29] ), .Z(\sub_109/carry[30] ) );
  XOR U885 ( .A(n1605), .B(\sub_109/carry[29] ), .Z(N32) );
  AND U886 ( .A(n523), .B(n524), .Z(terminate) );
  ANDN U887 ( .A(n525), .B(n526), .Z(n524) );
  ANDN U888 ( .A(n527), .B(n528), .Z(n525) );
  ANDN U889 ( .A(n529), .B(n530), .Z(n523) );
  ANDN U890 ( .A(iter[2]), .B(n531), .Z(n529) );
  IV U891 ( .A(n532), .Z(n1528) );
  IV U892 ( .A(n533), .Z(n1529) );
  IV U893 ( .A(n534), .Z(n1530) );
  IV U894 ( .A(n535), .Z(n1531) );
  IV U895 ( .A(n536), .Z(n1532) );
  IV U896 ( .A(n537), .Z(n1533) );
  IV U897 ( .A(n538), .Z(n1534) );
  IV U898 ( .A(n539), .Z(n1535) );
  IV U899 ( .A(n540), .Z(n1536) );
  IV U900 ( .A(n541), .Z(n1537) );
  IV U901 ( .A(n542), .Z(n1538) );
  IV U902 ( .A(n543), .Z(n1539) );
  IV U903 ( .A(n544), .Z(n1540) );
  IV U904 ( .A(n545), .Z(n1541) );
  IV U905 ( .A(n546), .Z(n1542) );
  IV U906 ( .A(n547), .Z(n1543) );
  IV U907 ( .A(n548), .Z(n1544) );
  IV U908 ( .A(n549), .Z(n1545) );
  IV U909 ( .A(n550), .Z(n1546) );
  IV U910 ( .A(n551), .Z(n1547) );
  IV U911 ( .A(n553), .Z(n1548) );
  IV U912 ( .A(n554), .Z(n1549) );
  IV U913 ( .A(n555), .Z(n1550) );
  IV U914 ( .A(n556), .Z(n1551) );
  IV U915 ( .A(n557), .Z(n1552) );
  IV U916 ( .A(n558), .Z(n1553) );
  IV U917 ( .A(n559), .Z(n1554) );
  IV U918 ( .A(n560), .Z(n1555) );
  IV U919 ( .A(n561), .Z(n1556) );
  IV U920 ( .A(n562), .Z(n1557) );
  IV U921 ( .A(n563), .Z(n1559) );
  IV U922 ( .A(n564), .Z(n1560) );
  IV U923 ( .A(n565), .Z(n1561) );
  IV U924 ( .A(n566), .Z(n1562) );
  IV U925 ( .A(n567), .Z(n1563) );
  IV U926 ( .A(n568), .Z(n1564) );
  IV U927 ( .A(n569), .Z(n1565) );
  IV U928 ( .A(n570), .Z(n1566) );
  IV U929 ( .A(n571), .Z(n1567) );
  IV U930 ( .A(n572), .Z(n1568) );
  IV U931 ( .A(n573), .Z(n1569) );
  IV U932 ( .A(n574), .Z(n1570) );
  IV U933 ( .A(n575), .Z(n1571) );
  IV U934 ( .A(n576), .Z(n1572) );
  IV U935 ( .A(n577), .Z(n1573) );
  IV U936 ( .A(n578), .Z(n1574) );
  IV U937 ( .A(n579), .Z(n1575) );
  IV U938 ( .A(n580), .Z(n1576) );
  IV U939 ( .A(n581), .Z(n1577) );
  IV U940 ( .A(n582), .Z(n1578) );
  IV U941 ( .A(n584), .Z(n1579) );
  IV U942 ( .A(n585), .Z(n1580) );
  IV U943 ( .A(n586), .Z(n1581) );
  IV U944 ( .A(n587), .Z(n1582) );
  IV U945 ( .A(n588), .Z(n1583) );
  IV U946 ( .A(n589), .Z(n1584) );
  IV U947 ( .A(n590), .Z(n1585) );
  IV U948 ( .A(n591), .Z(n1586) );
  IV U949 ( .A(n592), .Z(n1587) );
  IV U950 ( .A(n593), .Z(n1588) );
  IV U951 ( .A(n594), .Z(n1589) );
  IV U952 ( .A(n595), .Z(n1590) );
  IV U953 ( .A(n596), .Z(n1591) );
  IV U954 ( .A(n597), .Z(n1592) );
  IV U955 ( .A(n598), .Z(n1593) );
  IV U956 ( .A(n599), .Z(n1594) );
  IV U957 ( .A(n600), .Z(n1595) );
  IV U958 ( .A(n601), .Z(n1596) );
  IV U959 ( .A(n602), .Z(n1597) );
  IV U960 ( .A(n603), .Z(n1599) );
  IV U961 ( .A(n604), .Z(n1601) );
  IV U962 ( .A(n605), .Z(n1602) );
  IV U963 ( .A(n606), .Z(n1603) );
  IV U964 ( .A(n607), .Z(n1604) );
  IV U965 ( .A(n608), .Z(n1605) );
  IV U966 ( .A(n609), .Z(n1606) );
  IV U967 ( .A(n610), .Z(n1607) );
  IV U968 ( .A(n611), .Z(n1608) );
  IV U969 ( .A(n612), .Z(n1609) );
  IV U970 ( .A(n613), .Z(n1610) );
  IV U971 ( .A(n614), .Z(n1611) );
  IV U972 ( .A(n615), .Z(n1613) );
  IV U973 ( .A(n616), .Z(n1614) );
  IV U974 ( .A(n617), .Z(n1615) );
  IV U975 ( .A(n618), .Z(n1616) );
  IV U976 ( .A(n619), .Z(n1617) );
  XNOR U977 ( .A(n528), .B(n620), .Z(n518) );
  NANDN U978 ( .B(iter[5]), .A(n621), .Z(n516) );
  NANDN U979 ( .B(n622), .A(\add_181/carry[5] ), .Z(n621) );
  MUX U980 ( .IN0(N103), .IN1(iter[1]), .SEL(n622), .F(n514) );
  MUX U981 ( .IN0(N104), .IN1(iter[2]), .SEL(n622), .F(n512) );
  MUX U982 ( .IN0(N105), .IN1(iter[3]), .SEL(n622), .F(n510) );
  MUX U983 ( .IN0(N106), .IN1(iter[4]), .SEL(n622), .F(n508) );
  MUX U984 ( .IN0(n623), .IN1(o[28]), .SEL(n622), .F(n506) );
  XOR U985 ( .A(o[28]), .B(n624), .Z(n623) );
  MUX U986 ( .IN0(n625), .IN1(o[0]), .SEL(n622), .F(n505) );
  XNOR U987 ( .A(n1600), .B(o[0]), .Z(n625) );
  MUX U988 ( .IN0(n626), .IN1(o[1]), .SEL(n622), .F(n504) );
  XOR U989 ( .A(o[1]), .B(n627), .Z(n626) );
  MUX U990 ( .IN0(n628), .IN1(o[2]), .SEL(n622), .F(n503) );
  XOR U991 ( .A(o[2]), .B(n629), .Z(n628) );
  MUX U992 ( .IN0(n630), .IN1(o[3]), .SEL(n622), .F(n502) );
  XOR U993 ( .A(o[3]), .B(n631), .Z(n630) );
  MUX U994 ( .IN0(n632), .IN1(o[4]), .SEL(n622), .F(n501) );
  XOR U995 ( .A(o[4]), .B(n633), .Z(n632) );
  MUX U996 ( .IN0(n634), .IN1(o[5]), .SEL(n622), .F(n500) );
  XOR U997 ( .A(o[5]), .B(n635), .Z(n634) );
  MUX U998 ( .IN0(n636), .IN1(o[6]), .SEL(n622), .F(n499) );
  XOR U999 ( .A(o[6]), .B(n637), .Z(n636) );
  MUX U1000 ( .IN0(n638), .IN1(o[7]), .SEL(n622), .F(n498) );
  XOR U1001 ( .A(o[7]), .B(n639), .Z(n638) );
  MUX U1002 ( .IN0(n640), .IN1(o[8]), .SEL(n622), .F(n497) );
  XOR U1003 ( .A(o[8]), .B(n641), .Z(n640) );
  MUX U1004 ( .IN0(n642), .IN1(o[9]), .SEL(n622), .F(n496) );
  XOR U1005 ( .A(o[9]), .B(n643), .Z(n642) );
  MUX U1006 ( .IN0(n644), .IN1(o[10]), .SEL(n622), .F(n495) );
  XOR U1007 ( .A(o[10]), .B(n645), .Z(n644) );
  MUX U1008 ( .IN0(n646), .IN1(o[11]), .SEL(n622), .F(n494) );
  XOR U1009 ( .A(o[11]), .B(n647), .Z(n646) );
  MUX U1010 ( .IN0(n648), .IN1(o[12]), .SEL(n622), .F(n493) );
  XOR U1011 ( .A(o[12]), .B(n649), .Z(n648) );
  MUX U1012 ( .IN0(n650), .IN1(o[13]), .SEL(n622), .F(n492) );
  XOR U1013 ( .A(o[13]), .B(n651), .Z(n650) );
  MUX U1014 ( .IN0(n652), .IN1(o[14]), .SEL(n622), .F(n491) );
  XOR U1015 ( .A(o[14]), .B(n653), .Z(n652) );
  MUX U1016 ( .IN0(n654), .IN1(o[15]), .SEL(n622), .F(n490) );
  XOR U1017 ( .A(o[15]), .B(n655), .Z(n654) );
  MUX U1018 ( .IN0(n656), .IN1(o[16]), .SEL(n622), .F(n489) );
  XOR U1019 ( .A(o[16]), .B(n657), .Z(n656) );
  MUX U1020 ( .IN0(n658), .IN1(o[17]), .SEL(n622), .F(n488) );
  XOR U1021 ( .A(o[17]), .B(n659), .Z(n658) );
  MUX U1022 ( .IN0(n660), .IN1(o[18]), .SEL(n622), .F(n487) );
  XOR U1023 ( .A(o[18]), .B(n661), .Z(n660) );
  MUX U1024 ( .IN0(n662), .IN1(o[19]), .SEL(n622), .F(n486) );
  XOR U1025 ( .A(o[19]), .B(n663), .Z(n662) );
  MUX U1026 ( .IN0(n664), .IN1(o[20]), .SEL(n622), .F(n485) );
  XOR U1027 ( .A(o[20]), .B(n665), .Z(n664) );
  MUX U1028 ( .IN0(n666), .IN1(o[21]), .SEL(n622), .F(n484) );
  XOR U1029 ( .A(o[21]), .B(n667), .Z(n666) );
  MUX U1030 ( .IN0(n668), .IN1(o[22]), .SEL(n622), .F(n483) );
  XOR U1031 ( .A(o[22]), .B(n669), .Z(n668) );
  MUX U1032 ( .IN0(n670), .IN1(o[23]), .SEL(n622), .F(n482) );
  XOR U1033 ( .A(o[23]), .B(n671), .Z(n670) );
  MUX U1034 ( .IN0(n672), .IN1(o[24]), .SEL(n622), .F(n481) );
  XOR U1035 ( .A(o[24]), .B(n673), .Z(n672) );
  MUX U1036 ( .IN0(n674), .IN1(o[25]), .SEL(n622), .F(n480) );
  XOR U1037 ( .A(o[25]), .B(n675), .Z(n674) );
  MUX U1038 ( .IN0(n676), .IN1(o[26]), .SEL(n622), .F(n479) );
  XOR U1039 ( .A(o[26]), .B(n677), .Z(n676) );
  MUX U1040 ( .IN0(n678), .IN1(o[27]), .SEL(n622), .F(n478) );
  XOR U1041 ( .A(o[27]), .B(n679), .Z(n678) );
  MUX U1042 ( .IN0(n680), .IN1(o[29]), .SEL(n622), .F(n477) );
  XOR U1043 ( .A(o[29]), .B(n681), .Z(n680) );
  MUX U1044 ( .IN0(n682), .IN1(o[30]), .SEL(n622), .F(n476) );
  XNOR U1045 ( .A(o[30]), .B(n683), .Z(n682) );
  IV U1046 ( .A(n684), .Z(n475) );
  MUX U1047 ( .IN0(n685), .IN1(n686), .SEL(n620), .F(n684) );
  XNOR U1048 ( .A(n687), .B(n688), .Z(n686) );
  XOR U1049 ( .A(n689), .B(n690), .Z(n688) );
  XNOR U1050 ( .A(n685), .B(n691), .Z(n687) );
  ANDN U1051 ( .A(n692), .B(n683), .Z(n691) );
  XNOR U1052 ( .A(n690), .B(n689), .Z(n683) );
  NOR U1053 ( .A(o[31]), .B(\sub_109/carry[30] ), .Z(n689) );
  IV U1054 ( .A(n693), .Z(n690) );
  XNOR U1055 ( .A(o[30]), .B(n693), .Z(n692) );
  XOR U1056 ( .A(n694), .B(n695), .Z(n681) );
  MUX U1057 ( .IN0(n608), .IN1(N32), .SEL(n685), .F(n695) );
  NOR U1058 ( .A(n1618), .B(iter[0]), .Z(n608) );
  IV U1059 ( .A(n696), .Z(n1618) );
  XOR U1060 ( .A(n697), .B(n698), .Z(n624) );
  MUX U1061 ( .IN0(n696), .IN1(N31), .SEL(n685), .F(n698) );
  AND U1062 ( .A(n699), .B(n700), .Z(n696) );
  XOR U1063 ( .A(n701), .B(n702), .Z(n679) );
  MUX U1064 ( .IN0(n601), .IN1(N30), .SEL(n685), .F(n702) );
  NAND U1065 ( .A(n703), .B(n704), .Z(n601) );
  NAND U1066 ( .A(n705), .B(n699), .Z(n704) );
  NOR U1067 ( .A(n526), .B(n706), .Z(n705) );
  NAND U1068 ( .A(n707), .B(n699), .Z(n703) );
  ANDN U1069 ( .A(n700), .B(n528), .Z(n707) );
  XOR U1070 ( .A(n708), .B(n709), .Z(n677) );
  MUX U1071 ( .IN0(n615), .IN1(N29), .SEL(n685), .F(n709) );
  NANDN U1072 ( .B(n710), .A(n711), .Z(n615) );
  XOR U1073 ( .A(n712), .B(n713), .Z(n675) );
  MUX U1074 ( .IN0(n602), .IN1(N28), .SEL(n685), .F(n713) );
  NAND U1075 ( .A(n714), .B(n711), .Z(n602) );
  XOR U1076 ( .A(n715), .B(n716), .Z(n673) );
  MUX U1077 ( .IN0(n616), .IN1(N27), .SEL(n685), .F(n716) );
  NANDN U1078 ( .B(n717), .A(n718), .Z(n616) );
  XOR U1079 ( .A(n719), .B(n720), .Z(n671) );
  MUX U1080 ( .IN0(n609), .IN1(N26), .SEL(n685), .F(n720) );
  NAND U1081 ( .A(n718), .B(n721), .Z(n609) );
  ANDN U1082 ( .A(n722), .B(n717), .Z(n721) );
  AND U1083 ( .A(n723), .B(n724), .Z(n717) );
  ANDN U1084 ( .A(n526), .B(n725), .Z(n723) );
  NAND U1085 ( .A(n726), .B(n699), .Z(n722) );
  ANDN U1086 ( .A(n528), .B(n725), .Z(n726) );
  ANDN U1087 ( .A(n711), .B(n710), .Z(n718) );
  ANDN U1088 ( .A(n727), .B(n728), .Z(n710) );
  ANDN U1089 ( .A(n725), .B(n528), .Z(n727) );
  NAND U1090 ( .A(n724), .B(n729), .Z(n711) );
  ANDN U1091 ( .A(n725), .B(n526), .Z(n729) );
  XOR U1092 ( .A(n730), .B(n731), .Z(n669) );
  MUX U1093 ( .IN0(n732), .IN1(N25), .SEL(n685), .F(n731) );
  IV U1094 ( .A(n1598), .Z(n732) );
  ANDN U1095 ( .A(n733), .B(n734), .Z(n1598) );
  ANDN U1096 ( .A(n714), .B(n735), .Z(n733) );
  NANDN U1097 ( .B(n736), .A(n724), .Z(n714) );
  XOR U1098 ( .A(n737), .B(n738), .Z(n667) );
  MUX U1099 ( .IN0(n598), .IN1(N24), .SEL(n685), .F(n738) );
  NAND U1100 ( .A(n739), .B(n740), .Z(n598) );
  ANDN U1101 ( .A(n741), .B(n734), .Z(n740) );
  NAND U1102 ( .A(n742), .B(n700), .Z(n741) );
  NOR U1103 ( .A(n531), .B(n743), .Z(n742) );
  XOR U1104 ( .A(n744), .B(n745), .Z(n665) );
  MUX U1105 ( .IN0(n746), .IN1(N23), .SEL(n685), .F(n745) );
  IV U1106 ( .A(n1612), .Z(n746) );
  ANDN U1107 ( .A(n747), .B(n734), .Z(n1612) );
  ANDN U1108 ( .A(n748), .B(n735), .Z(n747) );
  NOR U1109 ( .A(n728), .B(n749), .Z(n735) );
  IV U1110 ( .A(n724), .Z(n728) );
  XOR U1111 ( .A(n750), .B(n751), .Z(n663) );
  MUX U1112 ( .IN0(n599), .IN1(N22), .SEL(n685), .F(n751) );
  NAND U1113 ( .A(n752), .B(n753), .Z(n599) );
  AND U1114 ( .A(n754), .B(n755), .Z(n753) );
  NANDN U1115 ( .B(n756), .A(n757), .Z(n755) );
  ANDN U1116 ( .A(n748), .B(n734), .Z(n754) );
  NAND U1117 ( .A(n758), .B(n759), .Z(n748) );
  ANDN U1118 ( .A(n526), .B(n531), .Z(n759) );
  AND U1119 ( .A(n760), .B(n761), .Z(n752) );
  NANDN U1120 ( .B(n762), .A(n699), .Z(n761) );
  NANDN U1121 ( .B(n763), .A(n699), .Z(n760) );
  XOR U1122 ( .A(n764), .B(n765), .Z(n661) );
  MUX U1123 ( .IN0(n617), .IN1(N21), .SEL(n685), .F(n765) );
  NAND U1124 ( .A(n766), .B(n739), .Z(n617) );
  AND U1125 ( .A(n767), .B(n768), .Z(n739) );
  NANDN U1126 ( .B(n528), .A(n724), .Z(n767) );
  XOR U1127 ( .A(n769), .B(n770), .Z(n659) );
  MUX U1128 ( .IN0(n610), .IN1(N20), .SEL(n685), .F(n770) );
  NAND U1129 ( .A(n766), .B(n771), .Z(n610) );
  OR U1130 ( .A(n772), .B(iter[0]), .Z(n771) );
  XOR U1131 ( .A(n773), .B(n774), .Z(n657) );
  MUX U1132 ( .IN0(n618), .IN1(N19), .SEL(n685), .F(n774) );
  NAND U1133 ( .A(n775), .B(n776), .Z(n618) );
  AND U1134 ( .A(n777), .B(n778), .Z(n776) );
  ANDN U1135 ( .A(n768), .B(n779), .Z(n778) );
  NANDN U1136 ( .B(n526), .A(n724), .Z(n768) );
  ANDN U1137 ( .A(n780), .B(n781), .Z(n775) );
  NAND U1138 ( .A(n782), .B(n699), .Z(n780) );
  AND U1139 ( .A(n531), .B(n530), .Z(n699) );
  ANDN U1140 ( .A(iter[0]), .B(n725), .Z(n782) );
  XOR U1141 ( .A(n783), .B(n784), .Z(n655) );
  MUX U1142 ( .IN0(n619), .IN1(N18), .SEL(n685), .F(n784) );
  NAND U1143 ( .A(n766), .B(n785), .Z(n619) );
  NOR U1144 ( .A(n781), .B(n786), .Z(n785) );
  NOR U1145 ( .A(n531), .B(n772), .Z(n781) );
  ANDN U1146 ( .A(n724), .B(n725), .Z(n734) );
  NOR U1147 ( .A(iter[4]), .B(iter[3]), .Z(n724) );
  NANDN U1148 ( .B(n531), .A(n758), .Z(n777) );
  XOR U1149 ( .A(n787), .B(n788), .Z(n653) );
  MUX U1150 ( .IN0(n611), .IN1(N17), .SEL(n685), .F(n788) );
  NAND U1151 ( .A(n789), .B(n790), .Z(n611) );
  AND U1152 ( .A(n791), .B(n792), .Z(n790) );
  XOR U1153 ( .A(n793), .B(n794), .Z(n651) );
  MUX U1154 ( .IN0(n603), .IN1(N16), .SEL(n685), .F(n794) );
  NAND U1155 ( .A(n795), .B(n796), .Z(n603) );
  AND U1156 ( .A(n797), .B(n798), .Z(n796) );
  ANDN U1157 ( .A(n799), .B(n758), .Z(n798) );
  ANDN U1158 ( .A(n800), .B(n786), .Z(n795) );
  XOR U1159 ( .A(n802), .B(n803), .Z(n649) );
  MUX U1160 ( .IN0(n604), .IN1(N15), .SEL(n685), .F(n803) );
  NAND U1161 ( .A(n804), .B(n805), .Z(n604) );
  ANDN U1162 ( .A(n806), .B(n779), .Z(n805) );
  AND U1163 ( .A(n799), .B(n807), .Z(n806) );
  AND U1164 ( .A(n791), .B(n808), .Z(n804) );
  NAND U1165 ( .A(iter[1]), .B(n809), .Z(n791) );
  XOR U1166 ( .A(n810), .B(n811), .Z(n647) );
  MUX U1167 ( .IN0(n597), .IN1(N14), .SEL(n685), .F(n811) );
  NAND U1168 ( .A(n812), .B(n813), .Z(n597) );
  AND U1169 ( .A(n799), .B(n814), .Z(n813) );
  ANDN U1170 ( .A(n807), .B(n815), .Z(n814) );
  NANDN U1171 ( .B(n816), .A(n801), .Z(n807) );
  AND U1172 ( .A(n797), .B(n817), .Z(n812) );
  NANDN U1173 ( .B(n818), .A(n757), .Z(n817) );
  XOR U1174 ( .A(n819), .B(n820), .Z(n645) );
  MUX U1175 ( .IN0(n612), .IN1(N13), .SEL(n685), .F(n820) );
  NAND U1176 ( .A(n789), .B(n821), .Z(n612) );
  ANDN U1177 ( .A(n792), .B(n822), .Z(n821) );
  NANDN U1178 ( .B(n528), .A(n530), .Z(n792) );
  AND U1179 ( .A(n823), .B(n799), .Z(n789) );
  NANDN U1180 ( .B(iter[1]), .A(n758), .Z(n823) );
  XOR U1181 ( .A(n824), .B(n825), .Z(n643) );
  MUX U1182 ( .IN0(n613), .IN1(N12), .SEL(n685), .F(n825) );
  NAND U1183 ( .A(n826), .B(n827), .Z(n613) );
  ANDN U1184 ( .A(n799), .B(n801), .Z(n827) );
  AND U1185 ( .A(n797), .B(n828), .Z(n826) );
  OR U1186 ( .A(n829), .B(iter[0]), .Z(n828) );
  NAND U1187 ( .A(iter[1]), .B(n530), .Z(n797) );
  XOR U1188 ( .A(n830), .B(n831), .Z(n641) );
  MUX U1189 ( .IN0(n605), .IN1(N11), .SEL(n685), .F(n831) );
  NAND U1190 ( .A(n832), .B(n833), .Z(n605) );
  ANDN U1191 ( .A(n834), .B(n822), .Z(n833) );
  AND U1192 ( .A(n835), .B(n836), .Z(n832) );
  XOR U1193 ( .A(n837), .B(n838), .Z(n639) );
  MUX U1194 ( .IN0(n595), .IN1(N10), .SEL(n685), .F(n838) );
  NAND U1195 ( .A(n839), .B(n840), .Z(n595) );
  AND U1196 ( .A(n834), .B(n841), .Z(n840) );
  ANDN U1197 ( .A(n842), .B(n843), .Z(n841) );
  ANDN U1198 ( .A(n799), .B(n844), .Z(n834) );
  ANDN U1199 ( .A(iter[4]), .B(n829), .Z(n844) );
  NANDN U1200 ( .B(iter[1]), .A(n531), .Z(n829) );
  ANDN U1201 ( .A(n845), .B(n779), .Z(n839) );
  AND U1202 ( .A(n528), .B(n758), .Z(n779) );
  ANDN U1203 ( .A(n846), .B(n822), .Z(n845) );
  AND U1204 ( .A(iter[4]), .B(n801), .Z(n822) );
  ANDN U1205 ( .A(n531), .B(iter[2]), .Z(n801) );
  OR U1206 ( .A(n818), .B(iter[0]), .Z(n846) );
  NANDN U1207 ( .B(iter[3]), .A(iter[4]), .Z(n818) );
  XOR U1208 ( .A(n847), .B(n848), .Z(n637) );
  MUX U1209 ( .IN0(n606), .IN1(N9), .SEL(n685), .F(n848) );
  NAND U1210 ( .A(n836), .B(n849), .Z(n606) );
  ANDN U1211 ( .A(n850), .B(n851), .Z(n849) );
  XOR U1212 ( .A(n852), .B(n853), .Z(n635) );
  MUX U1213 ( .IN0(n614), .IN1(N8), .SEL(n685), .F(n853) );
  NAND U1214 ( .A(n854), .B(n855), .Z(n614) );
  NOR U1215 ( .A(n786), .B(n843), .Z(n855) );
  AND U1216 ( .A(n528), .B(n530), .Z(n786) );
  ANDN U1217 ( .A(n856), .B(n851), .Z(n854) );
  NANDN U1218 ( .B(iter[0]), .A(n700), .Z(n856) );
  AND U1219 ( .A(n526), .B(n725), .Z(n700) );
  XOR U1220 ( .A(n857), .B(n858), .Z(n633) );
  MUX U1221 ( .IN0(n607), .IN1(N7), .SEL(n685), .F(n858) );
  NAND U1222 ( .A(n859), .B(n860), .Z(n607) );
  AND U1223 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U1224 ( .B(n528), .A(n863), .Z(n862) );
  AND U1225 ( .A(n850), .B(n864), .Z(n861) );
  OR U1226 ( .A(n762), .B(n865), .Z(n850) );
  NANDN U1227 ( .B(iter[0]), .A(iter[1]), .Z(n762) );
  ANDN U1228 ( .A(n836), .B(n866), .Z(n859) );
  ANDN U1229 ( .A(n808), .B(n867), .Z(n836) );
  XOR U1230 ( .A(n868), .B(n869), .Z(n631) );
  MUX U1231 ( .IN0(n594), .IN1(N6), .SEL(n685), .F(n869) );
  NAND U1232 ( .A(n870), .B(n871), .Z(n594) );
  AND U1233 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U1234 ( .B(n530), .A(n725), .Z(n873) );
  AND U1235 ( .A(n842), .B(n874), .Z(n872) );
  NANDN U1236 ( .B(n763), .A(n809), .Z(n874) );
  NANDN U1237 ( .B(iter[1]), .A(iter[0]), .Z(n763) );
  NANDN U1238 ( .B(n743), .A(iter[1]), .Z(n842) );
  NOR U1239 ( .A(n757), .B(n851), .Z(n870) );
  NAND U1240 ( .A(n799), .B(n875), .Z(n851) );
  NAND U1241 ( .A(iter[3]), .B(n530), .Z(n799) );
  ANDN U1242 ( .A(n725), .B(iter[0]), .Z(n757) );
  XOR U1243 ( .A(n876), .B(n877), .Z(n629) );
  MUX U1244 ( .IN0(n600), .IN1(N5), .SEL(n685), .F(n877) );
  NAND U1245 ( .A(n878), .B(n879), .Z(n600) );
  AND U1246 ( .A(n880), .B(n881), .Z(n879) );
  ANDN U1247 ( .A(n882), .B(n843), .Z(n881) );
  AND U1248 ( .A(iter[1]), .B(n758), .Z(n843) );
  AND U1249 ( .A(n883), .B(n875), .Z(n880) );
  AND U1250 ( .A(n884), .B(n885), .Z(n878) );
  AND U1251 ( .A(n864), .B(n886), .Z(n885) );
  NANDN U1252 ( .B(n526), .A(n887), .Z(n886) );
  ANDN U1253 ( .A(n530), .B(n528), .Z(n887) );
  AND U1254 ( .A(n888), .B(n889), .Z(n884) );
  NANDN U1255 ( .B(n528), .A(n758), .Z(n889) );
  OR U1256 ( .A(n736), .B(n725), .Z(n888) );
  NANDN U1257 ( .B(iter[0]), .A(n526), .Z(n736) );
  XOR U1258 ( .A(n890), .B(n891), .Z(n627) );
  MUX U1259 ( .IN0(n596), .IN1(N4), .SEL(n685), .F(n891) );
  NAND U1260 ( .A(n892), .B(n893), .Z(n596) );
  ANDN U1261 ( .A(n894), .B(n867), .Z(n893) );
  ANDN U1262 ( .A(iter[2]), .B(n772), .Z(n867) );
  ANDN U1263 ( .A(n882), .B(n815), .Z(n894) );
  ANDN U1264 ( .A(iter[2]), .B(n743), .Z(n815) );
  NANDN U1265 ( .B(iter[0]), .A(n530), .Z(n743) );
  NANDN U1266 ( .B(n706), .A(iter[4]), .Z(n882) );
  NANDN U1267 ( .B(iter[0]), .A(n725), .Z(n706) );
  AND U1268 ( .A(n895), .B(n896), .Z(n892) );
  ANDN U1269 ( .A(n897), .B(n866), .Z(n896) );
  OR U1270 ( .A(n749), .B(n865), .Z(n897) );
  IV U1271 ( .A(n758), .Z(n865) );
  ANDN U1272 ( .A(n530), .B(iter[2]), .Z(n758) );
  NANDN U1273 ( .B(n526), .A(iter[0]), .Z(n749) );
  MUX U1274 ( .IN0(n756), .IN1(n816), .SEL(iter[0]), .F(n895) );
  NANDN U1275 ( .B(n530), .A(n526), .Z(n816) );
  IV U1276 ( .A(n863), .Z(n756) );
  ANDN U1277 ( .A(o[0]), .B(n1600), .Z(n890) );
  AND U1278 ( .A(n898), .B(n899), .Z(n1600) );
  AND U1279 ( .A(n835), .B(n900), .Z(n899) );
  AND U1280 ( .A(n864), .B(n808), .Z(n900) );
  NAND U1281 ( .A(iter[0]), .B(n809), .Z(n808) );
  NAND U1282 ( .A(iter[4]), .B(n901), .Z(n864) );
  ANDN U1283 ( .A(n526), .B(iter[2]), .Z(n901) );
  OR U1284 ( .A(n772), .B(n528), .Z(n835) );
  NANDN U1285 ( .B(iter[1]), .A(n530), .Z(n772) );
  ANDN U1286 ( .A(n902), .B(n866), .Z(n898) );
  NAND U1287 ( .A(n883), .B(n875), .Z(n866) );
  NAND U1288 ( .A(iter[4]), .B(n531), .Z(n875) );
  NANDN U1289 ( .B(n531), .A(n809), .Z(n883) );
  AND U1290 ( .A(n530), .B(iter[2]), .Z(n809) );
  AND U1291 ( .A(n903), .B(n904), .Z(n902) );
  NANDN U1292 ( .B(n530), .A(n905), .Z(n904) );
  ANDN U1293 ( .A(n528), .B(n526), .Z(n905) );
  NANDN U1294 ( .B(n526), .A(n863), .Z(n903) );
  ANDN U1295 ( .A(n530), .B(n531), .Z(n863) );
  MUX U1296 ( .IN0(n906), .IN1(o[32]), .SEL(n622), .F(n474) );
  XOR U1297 ( .A(o[32]), .B(n907), .Z(n906) );
  IV U1298 ( .A(n908), .Z(n473) );
  MUX U1299 ( .IN0(n909), .IN1(n910), .SEL(n620), .F(n908) );
  XNOR U1300 ( .A(n909), .B(n911), .Z(n910) );
  IV U1301 ( .A(n912), .Z(n472) );
  MUX U1302 ( .IN0(n913), .IN1(n914), .SEL(n620), .F(n912) );
  XOR U1303 ( .A(n913), .B(n915), .Z(n914) );
  IV U1304 ( .A(n916), .Z(n471) );
  MUX U1305 ( .IN0(n917), .IN1(n918), .SEL(n620), .F(n916) );
  XOR U1306 ( .A(n917), .B(n919), .Z(n918) );
  IV U1307 ( .A(n920), .Z(n470) );
  MUX U1308 ( .IN0(n921), .IN1(n922), .SEL(n620), .F(n920) );
  XOR U1309 ( .A(n921), .B(n923), .Z(n922) );
  IV U1310 ( .A(n924), .Z(n469) );
  MUX U1311 ( .IN0(n925), .IN1(n926), .SEL(n620), .F(n924) );
  XOR U1312 ( .A(n925), .B(n927), .Z(n926) );
  IV U1313 ( .A(n928), .Z(n468) );
  MUX U1314 ( .IN0(n929), .IN1(n930), .SEL(n620), .F(n928) );
  XOR U1315 ( .A(n929), .B(n931), .Z(n930) );
  IV U1316 ( .A(n932), .Z(n467) );
  MUX U1317 ( .IN0(n933), .IN1(n934), .SEL(n620), .F(n932) );
  XOR U1318 ( .A(n933), .B(n935), .Z(n934) );
  IV U1319 ( .A(n936), .Z(n466) );
  MUX U1320 ( .IN0(n937), .IN1(n938), .SEL(n620), .F(n936) );
  XOR U1321 ( .A(n937), .B(n939), .Z(n938) );
  IV U1322 ( .A(n940), .Z(n465) );
  MUX U1323 ( .IN0(n941), .IN1(n942), .SEL(n620), .F(n940) );
  XOR U1324 ( .A(n941), .B(n943), .Z(n942) );
  IV U1325 ( .A(n944), .Z(n464) );
  MUX U1326 ( .IN0(n945), .IN1(n946), .SEL(n620), .F(n944) );
  XOR U1327 ( .A(n945), .B(n947), .Z(n946) );
  IV U1328 ( .A(n948), .Z(n463) );
  MUX U1329 ( .IN0(n949), .IN1(n950), .SEL(n620), .F(n948) );
  XOR U1330 ( .A(n949), .B(n951), .Z(n950) );
  MUX U1331 ( .IN0(n952), .IN1(o[44]), .SEL(n622), .F(n462) );
  XOR U1332 ( .A(o[44]), .B(n953), .Z(n952) );
  MUX U1333 ( .IN0(n954), .IN1(o[45]), .SEL(n622), .F(n461) );
  XOR U1334 ( .A(o[45]), .B(n955), .Z(n954) );
  MUX U1335 ( .IN0(n956), .IN1(o[46]), .SEL(n622), .F(n460) );
  XOR U1336 ( .A(o[46]), .B(n957), .Z(n956) );
  MUX U1337 ( .IN0(n958), .IN1(o[47]), .SEL(n622), .F(n459) );
  XOR U1338 ( .A(o[47]), .B(n959), .Z(n958) );
  MUX U1339 ( .IN0(n960), .IN1(o[48]), .SEL(n622), .F(n458) );
  XOR U1340 ( .A(o[48]), .B(n961), .Z(n960) );
  MUX U1341 ( .IN0(n962), .IN1(o[49]), .SEL(n622), .F(n457) );
  XOR U1342 ( .A(o[49]), .B(n963), .Z(n962) );
  MUX U1343 ( .IN0(n964), .IN1(o[50]), .SEL(n622), .F(n456) );
  XOR U1344 ( .A(o[50]), .B(n965), .Z(n964) );
  MUX U1345 ( .IN0(n966), .IN1(o[51]), .SEL(n622), .F(n455) );
  XOR U1346 ( .A(o[51]), .B(n967), .Z(n966) );
  MUX U1347 ( .IN0(n968), .IN1(o[52]), .SEL(n622), .F(n454) );
  XOR U1348 ( .A(o[52]), .B(n969), .Z(n968) );
  MUX U1349 ( .IN0(n970), .IN1(o[53]), .SEL(n622), .F(n453) );
  XOR U1350 ( .A(o[53]), .B(n971), .Z(n970) );
  MUX U1351 ( .IN0(n972), .IN1(o[54]), .SEL(n622), .F(n452) );
  XOR U1352 ( .A(o[54]), .B(n973), .Z(n972) );
  MUX U1353 ( .IN0(n974), .IN1(o[55]), .SEL(n622), .F(n451) );
  XOR U1354 ( .A(o[55]), .B(n975), .Z(n974) );
  MUX U1355 ( .IN0(n976), .IN1(o[56]), .SEL(n622), .F(n450) );
  XOR U1356 ( .A(o[56]), .B(n977), .Z(n976) );
  MUX U1357 ( .IN0(n978), .IN1(o[57]), .SEL(n622), .F(n449) );
  XOR U1358 ( .A(o[57]), .B(n979), .Z(n978) );
  MUX U1359 ( .IN0(n980), .IN1(o[58]), .SEL(n622), .F(n448) );
  XOR U1360 ( .A(o[58]), .B(n981), .Z(n980) );
  MUX U1361 ( .IN0(n982), .IN1(o[59]), .SEL(n622), .F(n447) );
  XOR U1362 ( .A(o[59]), .B(n983), .Z(n982) );
  MUX U1363 ( .IN0(n984), .IN1(o[60]), .SEL(n622), .F(n446) );
  XOR U1364 ( .A(o[60]), .B(n985), .Z(n984) );
  MUX U1365 ( .IN0(n986), .IN1(o[61]), .SEL(n622), .F(n445) );
  XOR U1366 ( .A(o[61]), .B(n987), .Z(n986) );
  IV U1367 ( .A(n988), .Z(n444) );
  MUX U1368 ( .IN0(n989), .IN1(n990), .SEL(n620), .F(n988) );
  XNOR U1369 ( .A(n989), .B(n991), .Z(n990) );
  MUX U1370 ( .IN0(n992), .IN1(o[63]), .SEL(n622), .F(n443) );
  XOR U1371 ( .A(n993), .B(n994), .Z(n992) );
  XOR U1372 ( .A(n995), .B(n996), .Z(n994) );
  MUX U1373 ( .IN0(N98), .IN1(n583), .SEL(n685), .F(n996) );
  AND U1374 ( .A(n997), .B(n998), .Z(n583) );
  XOR U1375 ( .A(o[63]), .B(n999), .Z(n993) );
  ANDN U1376 ( .A(n1000), .B(n991), .Z(n999) );
  XNOR U1377 ( .A(n995), .B(n1001), .Z(n991) );
  MUX U1378 ( .IN0(N97), .IN1(n575), .SEL(n685), .F(n1001) );
  ANDN U1379 ( .A(n998), .B(n1002), .Z(n575) );
  XNOR U1380 ( .A(n989), .B(n995), .Z(n1000) );
  XOR U1381 ( .A(n1003), .B(n1004), .Z(n987) );
  MUX U1382 ( .IN0(N96), .IN1(n587), .SEL(n685), .F(n1004) );
  AND U1383 ( .A(n1005), .B(n998), .Z(n587) );
  XOR U1384 ( .A(n1006), .B(n1007), .Z(n985) );
  MUX U1385 ( .IN0(N95), .IN1(n567), .SEL(n685), .F(n1007) );
  ANDN U1386 ( .A(n998), .B(n1008), .Z(n567) );
  XOR U1387 ( .A(n1009), .B(n1010), .Z(n983) );
  MUX U1388 ( .IN0(N94), .IN1(n579), .SEL(n685), .F(n1010) );
  AND U1389 ( .A(n1011), .B(n998), .Z(n579) );
  XOR U1390 ( .A(n1012), .B(n1013), .Z(n981) );
  MUX U1391 ( .IN0(N93), .IN1(n571), .SEL(n685), .F(n1013) );
  AND U1392 ( .A(n1014), .B(n998), .Z(n571) );
  XOR U1393 ( .A(n1015), .B(n1016), .Z(n979) );
  MUX U1394 ( .IN0(N92), .IN1(n592), .SEL(n685), .F(n1016) );
  AND U1395 ( .A(n1017), .B(n998), .Z(n592) );
  XOR U1396 ( .A(n1018), .B(n1019), .Z(n977) );
  MUX U1397 ( .IN0(N91), .IN1(n564), .SEL(n685), .F(n1019) );
  AND U1398 ( .A(n1020), .B(n998), .Z(n564) );
  XOR U1399 ( .A(n1021), .B(n1022), .Z(n975) );
  MUX U1400 ( .IN0(N90), .IN1(n584), .SEL(n685), .F(n1022) );
  AND U1401 ( .A(n1023), .B(n998), .Z(n584) );
  XOR U1402 ( .A(n1024), .B(n1025), .Z(n973) );
  MUX U1403 ( .IN0(N89), .IN1(n576), .SEL(n685), .F(n1025) );
  ANDN U1404 ( .A(n998), .B(n1026), .Z(n576) );
  XOR U1405 ( .A(n1027), .B(n1028), .Z(n971) );
  MUX U1406 ( .IN0(N88), .IN1(n588), .SEL(n685), .F(n1028) );
  AND U1407 ( .A(n1029), .B(n998), .Z(n588) );
  XOR U1408 ( .A(n1030), .B(n1031), .Z(n969) );
  MUX U1409 ( .IN0(N87), .IN1(n568), .SEL(n685), .F(n1031) );
  ANDN U1410 ( .A(n998), .B(n1032), .Z(n568) );
  XOR U1411 ( .A(n1033), .B(n1034), .Z(n967) );
  MUX U1412 ( .IN0(N86), .IN1(n580), .SEL(n685), .F(n1034) );
  AND U1413 ( .A(n1035), .B(n998), .Z(n580) );
  XOR U1414 ( .A(n1036), .B(n1037), .Z(n965) );
  MUX U1415 ( .IN0(N85), .IN1(n572), .SEL(n685), .F(n1037) );
  AND U1416 ( .A(n1038), .B(n998), .Z(n572) );
  XOR U1417 ( .A(n1039), .B(n1040), .Z(n963) );
  MUX U1418 ( .IN0(N84), .IN1(n590), .SEL(n685), .F(n1040) );
  AND U1419 ( .A(n1041), .B(n998), .Z(n590) );
  XOR U1420 ( .A(n1042), .B(n1043), .Z(n961) );
  MUX U1421 ( .IN0(N83), .IN1(n563), .SEL(n685), .F(n1043) );
  AND U1422 ( .A(n1044), .B(n998), .Z(n563) );
  XOR U1423 ( .A(n1045), .B(n1046), .Z(n959) );
  MUX U1424 ( .IN0(N82), .IN1(n582), .SEL(n685), .F(n1046) );
  ANDN U1425 ( .A(n1047), .B(iter[5]), .Z(n582) );
  MUX U1426 ( .IN0(n997), .IN1(n1048), .SEL(n530), .F(n1047) );
  MUX U1427 ( .IN0(n1049), .IN1(n1050), .SEL(iter[3]), .F(n1048) );
  AND U1428 ( .A(n1051), .B(n531), .Z(n997) );
  XOR U1429 ( .A(n1052), .B(n1053), .Z(n957) );
  MUX U1430 ( .IN0(N81), .IN1(n574), .SEL(n685), .F(n1053) );
  NOR U1431 ( .A(iter[5]), .B(n1054), .Z(n574) );
  MUX U1432 ( .IN0(n1055), .IN1(n1002), .SEL(iter[4]), .F(n1054) );
  OR U1433 ( .A(n1056), .B(iter[3]), .Z(n1002) );
  MUX U1434 ( .IN0(n1057), .IN1(n1058), .SEL(n531), .F(n1055) );
  XOR U1435 ( .A(n1059), .B(n1060), .Z(n955) );
  MUX U1436 ( .IN0(N80), .IN1(n586), .SEL(n685), .F(n1060) );
  ANDN U1437 ( .A(n1061), .B(iter[5]), .Z(n586) );
  MUX U1438 ( .IN0(n1005), .IN1(n1062), .SEL(n530), .F(n1061) );
  MUX U1439 ( .IN0(n1063), .IN1(n1064), .SEL(iter[3]), .F(n1062) );
  AND U1440 ( .A(n1065), .B(n531), .Z(n1005) );
  XOR U1441 ( .A(n1066), .B(n1067), .Z(n953) );
  MUX U1442 ( .IN0(N79), .IN1(n566), .SEL(n685), .F(n1067) );
  NOR U1443 ( .A(iter[5]), .B(n1068), .Z(n566) );
  MUX U1444 ( .IN0(n1069), .IN1(n1008), .SEL(iter[4]), .F(n1068) );
  OR U1445 ( .A(n1070), .B(iter[3]), .Z(n1008) );
  MUX U1446 ( .IN0(n1071), .IN1(n1072), .SEL(n531), .F(n1069) );
  XOR U1447 ( .A(n1073), .B(n1074), .Z(n951) );
  MUX U1448 ( .IN0(N78), .IN1(n578), .SEL(n685), .F(n1074) );
  ANDN U1449 ( .A(n1075), .B(iter[5]), .Z(n578) );
  MUX U1450 ( .IN0(n1011), .IN1(n1076), .SEL(n530), .F(n1075) );
  MUX U1451 ( .IN0(n1077), .IN1(n1078), .SEL(iter[3]), .F(n1076) );
  AND U1452 ( .A(n1079), .B(n531), .Z(n1011) );
  XOR U1453 ( .A(n1080), .B(n1081), .Z(n947) );
  MUX U1454 ( .IN0(N77), .IN1(n570), .SEL(n685), .F(n1081) );
  ANDN U1455 ( .A(n1082), .B(iter[5]), .Z(n570) );
  MUX U1456 ( .IN0(n1014), .IN1(n1083), .SEL(n530), .F(n1082) );
  MUX U1457 ( .IN0(n1084), .IN1(n1085), .SEL(iter[3]), .F(n1083) );
  AND U1458 ( .A(n1086), .B(n531), .Z(n1014) );
  XOR U1459 ( .A(n1087), .B(n1088), .Z(n943) );
  MUX U1460 ( .IN0(N76), .IN1(n593), .SEL(n685), .F(n1088) );
  ANDN U1461 ( .A(n1089), .B(iter[5]), .Z(n593) );
  MUX U1462 ( .IN0(n1017), .IN1(n1090), .SEL(n530), .F(n1089) );
  MUX U1463 ( .IN0(n1091), .IN1(n1092), .SEL(iter[3]), .F(n1090) );
  ANDN U1464 ( .A(n1093), .B(iter[3]), .Z(n1017) );
  XOR U1465 ( .A(n1094), .B(n1095), .Z(n939) );
  MUX U1466 ( .IN0(N75), .IN1(n565), .SEL(n685), .F(n1095) );
  ANDN U1467 ( .A(n1096), .B(iter[5]), .Z(n565) );
  MUX U1468 ( .IN0(n1020), .IN1(n1097), .SEL(n530), .F(n1096) );
  MUX U1469 ( .IN0(n1098), .IN1(n1099), .SEL(iter[3]), .F(n1097) );
  ANDN U1470 ( .A(n1100), .B(iter[3]), .Z(n1020) );
  XOR U1471 ( .A(n1101), .B(n1102), .Z(n935) );
  MUX U1472 ( .IN0(N74), .IN1(n585), .SEL(n685), .F(n1102) );
  ANDN U1473 ( .A(n1103), .B(iter[5]), .Z(n585) );
  MUX U1474 ( .IN0(n1023), .IN1(n1104), .SEL(n530), .F(n1103) );
  MUX U1475 ( .IN0(n1105), .IN1(n1049), .SEL(iter[3]), .F(n1104) );
  MUX U1476 ( .IN0(n1106), .IN1(n1107), .SEL(n725), .F(n1049) );
  MUX U1477 ( .IN0(n1108), .IN1(n1109), .SEL(n725), .F(n1105) );
  MUX U1478 ( .IN0(n1050), .IN1(n1051), .SEL(iter[3]), .F(n1023) );
  AND U1479 ( .A(n1110), .B(n725), .Z(n1051) );
  MUX U1480 ( .IN0(n1111), .IN1(n1112), .SEL(n725), .F(n1050) );
  XOR U1481 ( .A(n1113), .B(n1114), .Z(n931) );
  MUX U1482 ( .IN0(N73), .IN1(n577), .SEL(n685), .F(n1114) );
  NOR U1483 ( .A(iter[5]), .B(n1115), .Z(n577) );
  MUX U1484 ( .IN0(n1026), .IN1(n1116), .SEL(n530), .F(n1115) );
  MUX U1485 ( .IN0(n1117), .IN1(n1058), .SEL(iter[3]), .F(n1116) );
  IV U1486 ( .A(n1118), .Z(n1058) );
  MUX U1487 ( .IN0(n1119), .IN1(n1120), .SEL(iter[2]), .F(n1118) );
  MUX U1488 ( .IN0(n1121), .IN1(n1122), .SEL(n725), .F(n1117) );
  MUX U1489 ( .IN0(n1057), .IN1(n1056), .SEL(iter[3]), .F(n1026) );
  NANDN U1490 ( .B(iter[2]), .A(n1123), .Z(n1056) );
  IV U1491 ( .A(n1124), .Z(n1057) );
  MUX U1492 ( .IN0(n1125), .IN1(n1126), .SEL(iter[2]), .F(n1124) );
  XOR U1493 ( .A(n1127), .B(n1128), .Z(n927) );
  MUX U1494 ( .IN0(N72), .IN1(n589), .SEL(n685), .F(n1128) );
  ANDN U1495 ( .A(n1129), .B(iter[5]), .Z(n589) );
  MUX U1496 ( .IN0(n1029), .IN1(n1130), .SEL(n530), .F(n1129) );
  MUX U1497 ( .IN0(n1131), .IN1(n1063), .SEL(iter[3]), .F(n1130) );
  MUX U1498 ( .IN0(n1132), .IN1(n1133), .SEL(n725), .F(n1063) );
  MUX U1499 ( .IN0(n1134), .IN1(n1135), .SEL(n725), .F(n1131) );
  MUX U1500 ( .IN0(n1064), .IN1(n1065), .SEL(iter[3]), .F(n1029) );
  ANDN U1501 ( .A(n1136), .B(iter[2]), .Z(n1065) );
  MUX U1502 ( .IN0(n1137), .IN1(n1138), .SEL(n725), .F(n1064) );
  XOR U1503 ( .A(n1139), .B(n1140), .Z(n923) );
  MUX U1504 ( .IN0(N71), .IN1(n569), .SEL(n685), .F(n1140) );
  NOR U1505 ( .A(iter[5]), .B(n1141), .Z(n569) );
  MUX U1506 ( .IN0(n1032), .IN1(n1142), .SEL(n530), .F(n1141) );
  MUX U1507 ( .IN0(n1143), .IN1(n1072), .SEL(iter[3]), .F(n1142) );
  IV U1508 ( .A(n1144), .Z(n1072) );
  MUX U1509 ( .IN0(n1145), .IN1(n1146), .SEL(iter[2]), .F(n1144) );
  MUX U1510 ( .IN0(n1147), .IN1(n1148), .SEL(n725), .F(n1143) );
  MUX U1511 ( .IN0(n1071), .IN1(n1070), .SEL(iter[3]), .F(n1032) );
  NANDN U1512 ( .B(iter[2]), .A(n1149), .Z(n1070) );
  IV U1513 ( .A(n1150), .Z(n1071) );
  MUX U1514 ( .IN0(n1151), .IN1(n1152), .SEL(iter[2]), .F(n1150) );
  XOR U1515 ( .A(n1153), .B(n1154), .Z(n919) );
  MUX U1516 ( .IN0(N70), .IN1(n581), .SEL(n685), .F(n1154) );
  ANDN U1517 ( .A(n1155), .B(iter[5]), .Z(n581) );
  MUX U1518 ( .IN0(n1035), .IN1(n1156), .SEL(n530), .F(n1155) );
  MUX U1519 ( .IN0(n1157), .IN1(n1077), .SEL(iter[3]), .F(n1156) );
  MUX U1520 ( .IN0(n1107), .IN1(n1108), .SEL(n725), .F(n1077) );
  MUX U1521 ( .IN0(n1158), .IN1(n1159), .SEL(iter[1]), .F(n1108) );
  MUX U1522 ( .IN0(n1160), .IN1(n1161), .SEL(iter[1]), .F(n1107) );
  MUX U1523 ( .IN0(n1109), .IN1(n1162), .SEL(n725), .F(n1157) );
  MUX U1524 ( .IN0(n1163), .IN1(n1164), .SEL(iter[1]), .F(n1162) );
  IV U1525 ( .A(n1165), .Z(n1163) );
  MUX U1526 ( .IN0(n1166), .IN1(n1167), .SEL(n526), .F(n1109) );
  MUX U1527 ( .IN0(n1078), .IN1(n1079), .SEL(iter[3]), .F(n1035) );
  MUX U1528 ( .IN0(n1110), .IN1(n1111), .SEL(n725), .F(n1079) );
  MUX U1529 ( .IN0(n1168), .IN1(n1169), .SEL(iter[1]), .F(n1111) );
  ANDN U1530 ( .A(n1170), .B(iter[1]), .Z(n1110) );
  MUX U1531 ( .IN0(n1112), .IN1(n1106), .SEL(n725), .F(n1078) );
  MUX U1532 ( .IN0(n1171), .IN1(n1172), .SEL(iter[1]), .F(n1106) );
  MUX U1533 ( .IN0(n1173), .IN1(n1174), .SEL(iter[1]), .F(n1112) );
  XOR U1534 ( .A(n1175), .B(n1176), .Z(n915) );
  MUX U1535 ( .IN0(N69), .IN1(n573), .SEL(n685), .F(n1176) );
  ANDN U1536 ( .A(n1177), .B(iter[5]), .Z(n573) );
  MUX U1537 ( .IN0(n1038), .IN1(n1178), .SEL(n530), .F(n1177) );
  MUX U1538 ( .IN0(n1179), .IN1(n1084), .SEL(iter[3]), .F(n1178) );
  MUX U1539 ( .IN0(n1119), .IN1(n1180), .SEL(n725), .F(n1084) );
  IV U1540 ( .A(n1121), .Z(n1180) );
  MUX U1541 ( .IN0(n1181), .IN1(n1182), .SEL(iter[1]), .F(n1121) );
  IV U1542 ( .A(n1183), .Z(n1182) );
  MUX U1543 ( .IN0(n1184), .IN1(n1185), .SEL(iter[1]), .F(n1119) );
  IV U1544 ( .A(n1186), .Z(n1179) );
  MUX U1545 ( .IN0(n1187), .IN1(n1122), .SEL(iter[2]), .F(n1186) );
  MUX U1546 ( .IN0(n1188), .IN1(n1189), .SEL(iter[1]), .F(n1122) );
  MUX U1547 ( .IN0(n1190), .IN1(n1191), .SEL(n526), .F(n1187) );
  IV U1548 ( .A(n1192), .Z(n1191) );
  MUX U1549 ( .IN0(n1085), .IN1(n1086), .SEL(iter[3]), .F(n1038) );
  MUX U1550 ( .IN0(n1123), .IN1(n1126), .SEL(n725), .F(n1086) );
  MUX U1551 ( .IN0(n1193), .IN1(n1194), .SEL(iter[1]), .F(n1126) );
  AND U1552 ( .A(n1195), .B(n526), .Z(n1123) );
  MUX U1553 ( .IN0(n1125), .IN1(n1120), .SEL(n725), .F(n1085) );
  MUX U1554 ( .IN0(n1196), .IN1(n1197), .SEL(iter[1]), .F(n1120) );
  MUX U1555 ( .IN0(n1198), .IN1(n1199), .SEL(iter[1]), .F(n1125) );
  XOR U1556 ( .A(n1200), .B(n1201), .Z(n911) );
  MUX U1557 ( .IN0(N68), .IN1(n591), .SEL(n685), .F(n1201) );
  ANDN U1558 ( .A(n1202), .B(iter[5]), .Z(n591) );
  MUX U1559 ( .IN0(n1203), .IN1(n1041), .SEL(iter[4]), .F(n1202) );
  MUX U1560 ( .IN0(n1093), .IN1(n1092), .SEL(n531), .F(n1041) );
  MUX U1561 ( .IN0(n1132), .IN1(n1138), .SEL(iter[2]), .F(n1092) );
  MUX U1562 ( .IN0(n1172), .IN1(n1173), .SEL(iter[1]), .F(n1138) );
  MUX U1563 ( .IN0(o[88]), .IN1(o[87]), .SEL(n528), .F(n1173) );
  MUX U1564 ( .IN0(o[86]), .IN1(o[85]), .SEL(n528), .F(n1172) );
  MUX U1565 ( .IN0(n1161), .IN1(n1171), .SEL(iter[1]), .F(n1132) );
  MUX U1566 ( .IN0(o[84]), .IN1(o[83]), .SEL(n528), .F(n1171) );
  MUX U1567 ( .IN0(o[82]), .IN1(o[81]), .SEL(n528), .F(n1161) );
  MUX U1568 ( .IN0(n1136), .IN1(n1137), .SEL(n725), .F(n1093) );
  MUX U1569 ( .IN0(n1174), .IN1(n1168), .SEL(iter[1]), .F(n1137) );
  MUX U1570 ( .IN0(o[92]), .IN1(o[91]), .SEL(n528), .F(n1168) );
  MUX U1571 ( .IN0(o[90]), .IN1(o[89]), .SEL(n528), .F(n1174) );
  MUX U1572 ( .IN0(n1170), .IN1(n1169), .SEL(n526), .F(n1136) );
  MUX U1573 ( .IN0(o[93]), .IN1(o[94]), .SEL(iter[0]), .F(n1169) );
  AND U1574 ( .A(o[95]), .B(n528), .Z(n1170) );
  MUX U1575 ( .IN0(n1091), .IN1(n1204), .SEL(n531), .F(n1203) );
  MUX U1576 ( .IN0(n1205), .IN1(n1135), .SEL(iter[2]), .F(n1204) );
  MUX U1577 ( .IN0(n1164), .IN1(n1167), .SEL(iter[1]), .F(n1135) );
  MUX U1578 ( .IN0(o[72]), .IN1(o[71]), .SEL(n528), .F(n1167) );
  MUX U1579 ( .IN0(o[70]), .IN1(o[69]), .SEL(n528), .F(n1164) );
  IV U1580 ( .A(n1206), .Z(n1205) );
  MUX U1581 ( .IN0(n1207), .IN1(n1165), .SEL(iter[1]), .F(n1206) );
  MUX U1582 ( .IN0(n1208), .IN1(n1209), .SEL(iter[0]), .F(n1165) );
  MUX U1583 ( .IN0(n1210), .IN1(n1211), .SEL(n528), .F(n1207) );
  MUX U1584 ( .IN0(n1134), .IN1(n1133), .SEL(iter[2]), .F(n1091) );
  MUX U1585 ( .IN0(n1159), .IN1(n1160), .SEL(iter[1]), .F(n1133) );
  MUX U1586 ( .IN0(o[80]), .IN1(o[79]), .SEL(n528), .F(n1160) );
  MUX U1587 ( .IN0(o[78]), .IN1(o[77]), .SEL(n528), .F(n1159) );
  MUX U1588 ( .IN0(n1166), .IN1(n1158), .SEL(iter[1]), .F(n1134) );
  MUX U1589 ( .IN0(o[76]), .IN1(o[75]), .SEL(n528), .F(n1158) );
  MUX U1590 ( .IN0(o[74]), .IN1(o[73]), .SEL(n528), .F(n1166) );
  NANDN U1591 ( .B(n1558), .A(o[32]), .Z(n1200) );
  IV U1592 ( .A(n907), .Z(n1558) );
  AND U1593 ( .A(n1212), .B(n527), .Z(n907) );
  MUX U1594 ( .IN0(n1044), .IN1(n1213), .SEL(n530), .F(n1212) );
  MUX U1595 ( .IN0(n1214), .IN1(n1098), .SEL(iter[3]), .F(n1213) );
  MUX U1596 ( .IN0(n1145), .IN1(n1215), .SEL(n725), .F(n1098) );
  IV U1597 ( .A(n1147), .Z(n1215) );
  MUX U1598 ( .IN0(n1189), .IN1(n1181), .SEL(iter[1]), .F(n1147) );
  MUX U1599 ( .IN0(n1216), .IN1(n1217), .SEL(n528), .F(n1181) );
  MUX U1600 ( .IN0(n1218), .IN1(n1219), .SEL(n528), .F(n1189) );
  MUX U1601 ( .IN0(n1183), .IN1(n1184), .SEL(iter[1]), .F(n1145) );
  MUX U1602 ( .IN0(o[78]), .IN1(o[79]), .SEL(iter[0]), .F(n1184) );
  MUX U1603 ( .IN0(o[76]), .IN1(o[77]), .SEL(iter[0]), .F(n1183) );
  MUX U1604 ( .IN0(n1220), .IN1(n1221), .SEL(n725), .F(n1214) );
  MUX U1605 ( .IN0(n1222), .IN1(n1192), .SEL(iter[1]), .F(n1221) );
  MUX U1606 ( .IN0(o[67]), .IN1(o[66]), .SEL(n528), .F(n1192) );
  MUX U1607 ( .IN0(o[65]), .IN1(o[64]), .SEL(n528), .F(n1222) );
  IV U1608 ( .A(n1148), .Z(n1220) );
  MUX U1609 ( .IN0(n1190), .IN1(n1188), .SEL(iter[1]), .F(n1148) );
  MUX U1610 ( .IN0(n1223), .IN1(n1224), .SEL(n528), .F(n1188) );
  MUX U1611 ( .IN0(n1209), .IN1(n1225), .SEL(iter[0]), .F(n1190) );
  MUX U1612 ( .IN0(n1099), .IN1(n1100), .SEL(iter[3]), .F(n1044) );
  MUX U1613 ( .IN0(n1152), .IN1(n1149), .SEL(iter[2]), .F(n1100) );
  MUX U1614 ( .IN0(n1194), .IN1(n1195), .SEL(iter[1]), .F(n1149) );
  MUX U1615 ( .IN0(o[95]), .IN1(o[94]), .SEL(n528), .F(n1195) );
  MUX U1616 ( .IN0(o[92]), .IN1(o[93]), .SEL(iter[0]), .F(n1194) );
  MUX U1617 ( .IN0(n1199), .IN1(n1193), .SEL(iter[1]), .F(n1152) );
  MUX U1618 ( .IN0(o[91]), .IN1(o[90]), .SEL(n528), .F(n1193) );
  MUX U1619 ( .IN0(o[88]), .IN1(o[89]), .SEL(iter[0]), .F(n1199) );
  MUX U1620 ( .IN0(n1146), .IN1(n1151), .SEL(iter[2]), .F(n1099) );
  MUX U1621 ( .IN0(n1197), .IN1(n1198), .SEL(iter[1]), .F(n1151) );
  MUX U1622 ( .IN0(o[86]), .IN1(o[87]), .SEL(iter[0]), .F(n1198) );
  MUX U1623 ( .IN0(o[84]), .IN1(o[85]), .SEL(iter[0]), .F(n1197) );
  MUX U1624 ( .IN0(n1185), .IN1(n1196), .SEL(iter[1]), .F(n1146) );
  MUX U1625 ( .IN0(o[82]), .IN1(o[83]), .SEL(iter[0]), .F(n1196) );
  MUX U1626 ( .IN0(o[80]), .IN1(o[81]), .SEL(iter[0]), .F(n1185) );
  IV U1627 ( .A(o[62]), .Z(n989) );
  MUX U1628 ( .IN0(n1226), .IN1(o[64]), .SEL(n622), .F(n442) );
  XOR U1629 ( .A(o[64]), .B(n1227), .Z(n1226) );
  IV U1630 ( .A(n1228), .Z(n441) );
  MUX U1631 ( .IN0(n1211), .IN1(n1229), .SEL(n620), .F(n1228) );
  XNOR U1632 ( .A(n1211), .B(n1230), .Z(n1229) );
  IV U1633 ( .A(n1231), .Z(n440) );
  MUX U1634 ( .IN0(n1210), .IN1(n1232), .SEL(n620), .F(n1231) );
  XOR U1635 ( .A(n1210), .B(n1233), .Z(n1232) );
  IV U1636 ( .A(n1234), .Z(n439) );
  MUX U1637 ( .IN0(n1208), .IN1(n1235), .SEL(n620), .F(n1234) );
  XOR U1638 ( .A(n1208), .B(n1236), .Z(n1235) );
  IV U1639 ( .A(n1237), .Z(n438) );
  MUX U1640 ( .IN0(n1209), .IN1(n1238), .SEL(n620), .F(n1237) );
  XOR U1641 ( .A(n1209), .B(n1239), .Z(n1238) );
  IV U1642 ( .A(n1240), .Z(n437) );
  MUX U1643 ( .IN0(n1225), .IN1(n1241), .SEL(n620), .F(n1240) );
  XOR U1644 ( .A(n1225), .B(n1242), .Z(n1241) );
  IV U1645 ( .A(n1243), .Z(n436) );
  MUX U1646 ( .IN0(n1224), .IN1(n1244), .SEL(n620), .F(n1243) );
  XOR U1647 ( .A(n1224), .B(n1245), .Z(n1244) );
  IV U1648 ( .A(n1246), .Z(n435) );
  MUX U1649 ( .IN0(n1223), .IN1(n1247), .SEL(n620), .F(n1246) );
  XOR U1650 ( .A(n1223), .B(n1248), .Z(n1247) );
  IV U1651 ( .A(n1249), .Z(n434) );
  MUX U1652 ( .IN0(n1219), .IN1(n1250), .SEL(n620), .F(n1249) );
  XOR U1653 ( .A(n1219), .B(n1251), .Z(n1250) );
  IV U1654 ( .A(n1252), .Z(n433) );
  MUX U1655 ( .IN0(n1218), .IN1(n1253), .SEL(n620), .F(n1252) );
  XOR U1656 ( .A(n1218), .B(n1254), .Z(n1253) );
  IV U1657 ( .A(n1255), .Z(n432) );
  MUX U1658 ( .IN0(n1217), .IN1(n1256), .SEL(n620), .F(n1255) );
  XOR U1659 ( .A(n1217), .B(n1257), .Z(n1256) );
  IV U1660 ( .A(n1258), .Z(n431) );
  MUX U1661 ( .IN0(n1216), .IN1(n1259), .SEL(n620), .F(n1258) );
  XOR U1662 ( .A(n1216), .B(n1260), .Z(n1259) );
  MUX U1663 ( .IN0(n1261), .IN1(o[76]), .SEL(n622), .F(n430) );
  XOR U1664 ( .A(o[76]), .B(n1262), .Z(n1261) );
  MUX U1665 ( .IN0(n1263), .IN1(o[77]), .SEL(n622), .F(n429) );
  XOR U1666 ( .A(o[77]), .B(n1264), .Z(n1263) );
  MUX U1667 ( .IN0(n1265), .IN1(o[78]), .SEL(n622), .F(n428) );
  XOR U1668 ( .A(o[78]), .B(n1266), .Z(n1265) );
  MUX U1669 ( .IN0(n1267), .IN1(o[79]), .SEL(n622), .F(n427) );
  XOR U1670 ( .A(o[79]), .B(n1268), .Z(n1267) );
  MUX U1671 ( .IN0(n1269), .IN1(o[80]), .SEL(n622), .F(n426) );
  XOR U1672 ( .A(o[80]), .B(n1270), .Z(n1269) );
  MUX U1673 ( .IN0(n1271), .IN1(o[81]), .SEL(n622), .F(n425) );
  XOR U1674 ( .A(o[81]), .B(n1272), .Z(n1271) );
  MUX U1675 ( .IN0(n1273), .IN1(o[82]), .SEL(n622), .F(n424) );
  XOR U1676 ( .A(o[82]), .B(n1274), .Z(n1273) );
  MUX U1677 ( .IN0(n1275), .IN1(o[83]), .SEL(n622), .F(n423) );
  XOR U1678 ( .A(o[83]), .B(n1276), .Z(n1275) );
  MUX U1679 ( .IN0(n1277), .IN1(o[84]), .SEL(n622), .F(n422) );
  XOR U1680 ( .A(o[84]), .B(n1278), .Z(n1277) );
  MUX U1681 ( .IN0(n1279), .IN1(o[85]), .SEL(n622), .F(n421) );
  XOR U1682 ( .A(o[85]), .B(n1280), .Z(n1279) );
  MUX U1683 ( .IN0(n1281), .IN1(o[86]), .SEL(n622), .F(n420) );
  XOR U1684 ( .A(o[86]), .B(n1282), .Z(n1281) );
  MUX U1685 ( .IN0(n1283), .IN1(o[87]), .SEL(n622), .F(n419) );
  XOR U1686 ( .A(o[87]), .B(n1284), .Z(n1283) );
  MUX U1687 ( .IN0(n1285), .IN1(o[88]), .SEL(n622), .F(n418) );
  XOR U1688 ( .A(o[88]), .B(n1286), .Z(n1285) );
  MUX U1689 ( .IN0(n1287), .IN1(o[89]), .SEL(n622), .F(n417) );
  XOR U1690 ( .A(o[89]), .B(n1288), .Z(n1287) );
  MUX U1691 ( .IN0(n1289), .IN1(o[90]), .SEL(n622), .F(n416) );
  XOR U1692 ( .A(o[90]), .B(n1290), .Z(n1289) );
  MUX U1693 ( .IN0(n1291), .IN1(o[91]), .SEL(n622), .F(n415) );
  XOR U1694 ( .A(o[91]), .B(n1292), .Z(n1291) );
  MUX U1695 ( .IN0(o[92]), .IN1(n1293), .SEL(n620), .F(n414) );
  XOR U1696 ( .A(o[92]), .B(n1294), .Z(n1293) );
  MUX U1697 ( .IN0(o[93]), .IN1(n1295), .SEL(n620), .F(n413) );
  XOR U1698 ( .A(o[93]), .B(n1296), .Z(n1295) );
  IV U1699 ( .A(n1297), .Z(n412) );
  MUX U1700 ( .IN0(n1298), .IN1(n1299), .SEL(n622), .F(n1297) );
  IV U1701 ( .A(n620), .Z(n622) );
  XNOR U1702 ( .A(n1299), .B(n1300), .Z(n1298) );
  MUX U1703 ( .IN0(o[95]), .IN1(n1301), .SEL(n620), .F(n411) );
  ANDN U1704 ( .A(n1302), .B(iter[5]), .Z(n620) );
  NAND U1705 ( .A(n1303), .B(n1304), .Z(n1302) );
  ANDN U1706 ( .A(n1305), .B(n725), .Z(n1304) );
  ANDN U1707 ( .A(iter[0]), .B(n526), .Z(n1305) );
  ANDN U1708 ( .A(iter[3]), .B(n530), .Z(n1303) );
  XOR U1709 ( .A(n1306), .B(n1307), .Z(n1301) );
  XOR U1710 ( .A(n1308), .B(n1309), .Z(n1307) );
  MUX U1711 ( .IN0(n552), .IN1(N66), .SEL(n685), .F(n1309) );
  AND U1712 ( .A(n1310), .B(n998), .Z(n552) );
  XOR U1713 ( .A(o[95]), .B(n1311), .Z(n1306) );
  ANDN U1714 ( .A(n1312), .B(n1300), .Z(n1311) );
  XNOR U1715 ( .A(n1308), .B(n1313), .Z(n1300) );
  MUX U1716 ( .IN0(n544), .IN1(N65), .SEL(n685), .F(n1313) );
  ANDN U1717 ( .A(n998), .B(n1314), .Z(n544) );
  XNOR U1718 ( .A(n1299), .B(n1308), .Z(n1312) );
  XOR U1719 ( .A(n1315), .B(n1316), .Z(n1296) );
  MUX U1720 ( .IN0(n556), .IN1(N64), .SEL(n685), .F(n1316) );
  AND U1721 ( .A(n1317), .B(n998), .Z(n556) );
  XOR U1722 ( .A(n1318), .B(n1319), .Z(n1294) );
  MUX U1723 ( .IN0(n536), .IN1(N63), .SEL(n685), .F(n1319) );
  ANDN U1724 ( .A(n998), .B(n1320), .Z(n536) );
  XOR U1725 ( .A(n1321), .B(n1322), .Z(n1292) );
  MUX U1726 ( .IN0(n548), .IN1(N62), .SEL(n685), .F(n1322) );
  AND U1727 ( .A(n1323), .B(n998), .Z(n548) );
  XOR U1728 ( .A(n1324), .B(n1325), .Z(n1290) );
  MUX U1729 ( .IN0(n540), .IN1(N61), .SEL(n685), .F(n1325) );
  AND U1730 ( .A(n1326), .B(n998), .Z(n540) );
  XOR U1731 ( .A(n1327), .B(n1328), .Z(n1288) );
  MUX U1732 ( .IN0(n561), .IN1(N60), .SEL(n685), .F(n1328) );
  AND U1733 ( .A(n1329), .B(n998), .Z(n561) );
  XOR U1734 ( .A(n1330), .B(n1331), .Z(n1286) );
  MUX U1735 ( .IN0(n533), .IN1(N59), .SEL(n685), .F(n1331) );
  AND U1736 ( .A(n1332), .B(n998), .Z(n533) );
  XOR U1737 ( .A(n1333), .B(n1334), .Z(n1284) );
  MUX U1738 ( .IN0(n553), .IN1(N58), .SEL(n685), .F(n1334) );
  AND U1739 ( .A(n1335), .B(n998), .Z(n553) );
  XOR U1740 ( .A(n1336), .B(n1337), .Z(n1282) );
  MUX U1741 ( .IN0(n545), .IN1(N57), .SEL(n685), .F(n1337) );
  ANDN U1742 ( .A(n998), .B(n1338), .Z(n545) );
  XOR U1743 ( .A(n1339), .B(n1340), .Z(n1280) );
  MUX U1744 ( .IN0(n557), .IN1(N56), .SEL(n685), .F(n1340) );
  AND U1745 ( .A(n1341), .B(n998), .Z(n557) );
  XOR U1746 ( .A(n1342), .B(n1343), .Z(n1278) );
  MUX U1747 ( .IN0(n537), .IN1(N55), .SEL(n685), .F(n1343) );
  ANDN U1748 ( .A(n998), .B(n1344), .Z(n537) );
  XOR U1749 ( .A(n1345), .B(n1346), .Z(n1276) );
  MUX U1750 ( .IN0(n549), .IN1(N54), .SEL(n685), .F(n1346) );
  AND U1751 ( .A(n1347), .B(n998), .Z(n549) );
  XOR U1752 ( .A(n1348), .B(n1349), .Z(n1274) );
  MUX U1753 ( .IN0(n541), .IN1(N53), .SEL(n685), .F(n1349) );
  AND U1754 ( .A(n1350), .B(n998), .Z(n541) );
  XOR U1755 ( .A(n1351), .B(n1352), .Z(n1272) );
  MUX U1756 ( .IN0(n559), .IN1(N52), .SEL(n685), .F(n1352) );
  AND U1757 ( .A(n1353), .B(n998), .Z(n559) );
  XOR U1758 ( .A(n1354), .B(n1355), .Z(n1270) );
  MUX U1759 ( .IN0(n532), .IN1(N51), .SEL(n685), .F(n1355) );
  AND U1760 ( .A(n1356), .B(n998), .Z(n532) );
  AND U1761 ( .A(n530), .B(n527), .Z(n998) );
  XOR U1762 ( .A(n1357), .B(n1358), .Z(n1268) );
  MUX U1763 ( .IN0(n551), .IN1(N50), .SEL(n685), .F(n1358) );
  ANDN U1764 ( .A(n1359), .B(iter[5]), .Z(n551) );
  MUX U1765 ( .IN0(n1310), .IN1(n1360), .SEL(n530), .F(n1359) );
  MUX U1766 ( .IN0(n1361), .IN1(n1362), .SEL(iter[3]), .F(n1360) );
  AND U1767 ( .A(n1363), .B(n531), .Z(n1310) );
  XOR U1768 ( .A(n1364), .B(n1365), .Z(n1266) );
  MUX U1769 ( .IN0(n543), .IN1(N49), .SEL(n685), .F(n1365) );
  NOR U1770 ( .A(iter[5]), .B(n1366), .Z(n543) );
  MUX U1771 ( .IN0(n1367), .IN1(n1314), .SEL(iter[4]), .F(n1366) );
  OR U1772 ( .A(n1368), .B(iter[3]), .Z(n1314) );
  MUX U1773 ( .IN0(n1369), .IN1(n1370), .SEL(n531), .F(n1367) );
  XOR U1774 ( .A(n1371), .B(n1372), .Z(n1264) );
  MUX U1775 ( .IN0(n555), .IN1(N48), .SEL(n685), .F(n1372) );
  ANDN U1776 ( .A(n1373), .B(iter[5]), .Z(n555) );
  MUX U1777 ( .IN0(n1317), .IN1(n1374), .SEL(n530), .F(n1373) );
  MUX U1778 ( .IN0(n1375), .IN1(n1376), .SEL(iter[3]), .F(n1374) );
  AND U1779 ( .A(n1377), .B(n531), .Z(n1317) );
  XOR U1780 ( .A(n1378), .B(n1379), .Z(n1262) );
  MUX U1781 ( .IN0(n535), .IN1(N47), .SEL(n685), .F(n1379) );
  NOR U1782 ( .A(iter[5]), .B(n1380), .Z(n535) );
  MUX U1783 ( .IN0(n1381), .IN1(n1320), .SEL(iter[4]), .F(n1380) );
  OR U1784 ( .A(n1382), .B(iter[3]), .Z(n1320) );
  MUX U1785 ( .IN0(n1383), .IN1(n1384), .SEL(n531), .F(n1381) );
  IV U1786 ( .A(o[75]), .Z(n1216) );
  XOR U1787 ( .A(n1385), .B(n1386), .Z(n1260) );
  MUX U1788 ( .IN0(n547), .IN1(N46), .SEL(n685), .F(n1386) );
  ANDN U1789 ( .A(n1387), .B(iter[5]), .Z(n547) );
  MUX U1790 ( .IN0(n1323), .IN1(n1388), .SEL(n530), .F(n1387) );
  MUX U1791 ( .IN0(n1389), .IN1(n1390), .SEL(iter[3]), .F(n1388) );
  AND U1792 ( .A(n1391), .B(n531), .Z(n1323) );
  IV U1793 ( .A(o[74]), .Z(n1217) );
  XOR U1794 ( .A(n1392), .B(n1393), .Z(n1257) );
  MUX U1795 ( .IN0(n539), .IN1(N45), .SEL(n685), .F(n1393) );
  ANDN U1796 ( .A(n1394), .B(iter[5]), .Z(n539) );
  MUX U1797 ( .IN0(n1326), .IN1(n1395), .SEL(n530), .F(n1394) );
  MUX U1798 ( .IN0(n1396), .IN1(n1397), .SEL(iter[3]), .F(n1395) );
  AND U1799 ( .A(n1398), .B(n531), .Z(n1326) );
  IV U1800 ( .A(o[73]), .Z(n1218) );
  XOR U1801 ( .A(n1399), .B(n1400), .Z(n1254) );
  MUX U1802 ( .IN0(n562), .IN1(N44), .SEL(n685), .F(n1400) );
  ANDN U1803 ( .A(n1401), .B(iter[5]), .Z(n562) );
  MUX U1804 ( .IN0(n1329), .IN1(n1402), .SEL(n530), .F(n1401) );
  MUX U1805 ( .IN0(n1403), .IN1(n1404), .SEL(iter[3]), .F(n1402) );
  ANDN U1806 ( .A(n1405), .B(iter[3]), .Z(n1329) );
  IV U1807 ( .A(o[72]), .Z(n1219) );
  XOR U1808 ( .A(n1406), .B(n1407), .Z(n1251) );
  MUX U1809 ( .IN0(n534), .IN1(N43), .SEL(n685), .F(n1407) );
  ANDN U1810 ( .A(n1408), .B(iter[5]), .Z(n534) );
  MUX U1811 ( .IN0(n1332), .IN1(n1409), .SEL(n530), .F(n1408) );
  MUX U1812 ( .IN0(n1410), .IN1(n1411), .SEL(iter[3]), .F(n1409) );
  ANDN U1813 ( .A(n1412), .B(iter[3]), .Z(n1332) );
  IV U1814 ( .A(o[71]), .Z(n1223) );
  XOR U1815 ( .A(n1413), .B(n1414), .Z(n1248) );
  MUX U1816 ( .IN0(n554), .IN1(N42), .SEL(n685), .F(n1414) );
  ANDN U1817 ( .A(n1415), .B(iter[5]), .Z(n554) );
  MUX U1818 ( .IN0(n1335), .IN1(n1416), .SEL(n530), .F(n1415) );
  MUX U1819 ( .IN0(n1417), .IN1(n1361), .SEL(iter[3]), .F(n1416) );
  MUX U1820 ( .IN0(n1418), .IN1(n1419), .SEL(n725), .F(n1361) );
  MUX U1821 ( .IN0(n1420), .IN1(n1421), .SEL(n725), .F(n1417) );
  MUX U1822 ( .IN0(n1362), .IN1(n1363), .SEL(iter[3]), .F(n1335) );
  AND U1823 ( .A(n1422), .B(n725), .Z(n1363) );
  MUX U1824 ( .IN0(n1423), .IN1(n1424), .SEL(n725), .F(n1362) );
  IV U1825 ( .A(o[70]), .Z(n1224) );
  XOR U1826 ( .A(n1425), .B(n1426), .Z(n1245) );
  MUX U1827 ( .IN0(n546), .IN1(N41), .SEL(n685), .F(n1426) );
  NOR U1828 ( .A(iter[5]), .B(n1427), .Z(n546) );
  MUX U1829 ( .IN0(n1338), .IN1(n1428), .SEL(n530), .F(n1427) );
  MUX U1830 ( .IN0(n1429), .IN1(n1370), .SEL(iter[3]), .F(n1428) );
  IV U1831 ( .A(n1430), .Z(n1370) );
  MUX U1832 ( .IN0(n1431), .IN1(n1432), .SEL(iter[2]), .F(n1430) );
  MUX U1833 ( .IN0(n1433), .IN1(n1434), .SEL(n725), .F(n1429) );
  MUX U1834 ( .IN0(n1369), .IN1(n1368), .SEL(iter[3]), .F(n1338) );
  NANDN U1835 ( .B(iter[2]), .A(n1435), .Z(n1368) );
  IV U1836 ( .A(n1436), .Z(n1369) );
  MUX U1837 ( .IN0(n1437), .IN1(n1438), .SEL(iter[2]), .F(n1436) );
  IV U1838 ( .A(o[69]), .Z(n1225) );
  XOR U1839 ( .A(n1439), .B(n1440), .Z(n1242) );
  MUX U1840 ( .IN0(n558), .IN1(N40), .SEL(n685), .F(n1440) );
  ANDN U1841 ( .A(n1441), .B(iter[5]), .Z(n558) );
  MUX U1842 ( .IN0(n1341), .IN1(n1442), .SEL(n530), .F(n1441) );
  MUX U1843 ( .IN0(n1443), .IN1(n1375), .SEL(iter[3]), .F(n1442) );
  MUX U1844 ( .IN0(n1444), .IN1(n1445), .SEL(n725), .F(n1375) );
  MUX U1845 ( .IN0(n1446), .IN1(n1447), .SEL(n725), .F(n1443) );
  MUX U1846 ( .IN0(n1376), .IN1(n1377), .SEL(iter[3]), .F(n1341) );
  ANDN U1847 ( .A(n1448), .B(iter[2]), .Z(n1377) );
  MUX U1848 ( .IN0(n1449), .IN1(n1450), .SEL(n725), .F(n1376) );
  IV U1849 ( .A(o[68]), .Z(n1209) );
  XOR U1850 ( .A(n1451), .B(n1452), .Z(n1239) );
  MUX U1851 ( .IN0(n538), .IN1(N39), .SEL(n685), .F(n1452) );
  NOR U1852 ( .A(iter[5]), .B(n1453), .Z(n538) );
  MUX U1853 ( .IN0(n1344), .IN1(n1454), .SEL(n530), .F(n1453) );
  MUX U1854 ( .IN0(n1455), .IN1(n1384), .SEL(iter[3]), .F(n1454) );
  IV U1855 ( .A(n1456), .Z(n1384) );
  MUX U1856 ( .IN0(n1457), .IN1(n1458), .SEL(iter[2]), .F(n1456) );
  MUX U1857 ( .IN0(n1459), .IN1(n1460), .SEL(n725), .F(n1455) );
  MUX U1858 ( .IN0(n1383), .IN1(n1382), .SEL(iter[3]), .F(n1344) );
  NANDN U1859 ( .B(iter[2]), .A(n1461), .Z(n1382) );
  IV U1860 ( .A(n1462), .Z(n1383) );
  MUX U1861 ( .IN0(n1463), .IN1(n1464), .SEL(iter[2]), .F(n1462) );
  IV U1862 ( .A(o[67]), .Z(n1208) );
  XOR U1863 ( .A(n1465), .B(n1466), .Z(n1236) );
  MUX U1864 ( .IN0(n550), .IN1(N38), .SEL(n685), .F(n1466) );
  ANDN U1865 ( .A(n1467), .B(iter[5]), .Z(n550) );
  MUX U1866 ( .IN0(n1347), .IN1(n1468), .SEL(n530), .F(n1467) );
  MUX U1867 ( .IN0(n1469), .IN1(n1389), .SEL(iter[3]), .F(n1468) );
  MUX U1868 ( .IN0(n1419), .IN1(n1420), .SEL(n725), .F(n1389) );
  MUX U1869 ( .IN0(n1470), .IN1(n1471), .SEL(iter[1]), .F(n1420) );
  MUX U1870 ( .IN0(n1472), .IN1(n1473), .SEL(iter[1]), .F(n1419) );
  MUX U1871 ( .IN0(n1421), .IN1(n1474), .SEL(n725), .F(n1469) );
  MUX U1872 ( .IN0(n1475), .IN1(n1476), .SEL(iter[1]), .F(n1474) );
  IV U1873 ( .A(n1477), .Z(n1475) );
  MUX U1874 ( .IN0(n1478), .IN1(n1479), .SEL(n526), .F(n1421) );
  MUX U1875 ( .IN0(n1390), .IN1(n1391), .SEL(iter[3]), .F(n1347) );
  MUX U1876 ( .IN0(n1422), .IN1(n1423), .SEL(n725), .F(n1391) );
  MUX U1877 ( .IN0(n1480), .IN1(n1481), .SEL(iter[1]), .F(n1423) );
  ANDN U1878 ( .A(n1482), .B(iter[1]), .Z(n1422) );
  MUX U1879 ( .IN0(n1424), .IN1(n1418), .SEL(n725), .F(n1390) );
  MUX U1880 ( .IN0(n1483), .IN1(n1484), .SEL(iter[1]), .F(n1418) );
  MUX U1881 ( .IN0(n1485), .IN1(n1486), .SEL(iter[1]), .F(n1424) );
  IV U1882 ( .A(o[66]), .Z(n1210) );
  XOR U1883 ( .A(n1487), .B(n1488), .Z(n1233) );
  MUX U1884 ( .IN0(n542), .IN1(N37), .SEL(n685), .F(n1488) );
  ANDN U1885 ( .A(n1489), .B(iter[5]), .Z(n542) );
  MUX U1886 ( .IN0(n1350), .IN1(n1490), .SEL(n530), .F(n1489) );
  MUX U1887 ( .IN0(n1491), .IN1(n1396), .SEL(iter[3]), .F(n1490) );
  MUX U1888 ( .IN0(n1431), .IN1(n1492), .SEL(n725), .F(n1396) );
  IV U1889 ( .A(n1433), .Z(n1492) );
  MUX U1890 ( .IN0(n1493), .IN1(n1494), .SEL(iter[1]), .F(n1433) );
  IV U1891 ( .A(n1495), .Z(n1494) );
  MUX U1892 ( .IN0(n1496), .IN1(n1497), .SEL(iter[1]), .F(n1431) );
  IV U1893 ( .A(n1498), .Z(n1491) );
  MUX U1894 ( .IN0(n1499), .IN1(n1434), .SEL(iter[2]), .F(n1498) );
  MUX U1895 ( .IN0(n1500), .IN1(n1501), .SEL(iter[1]), .F(n1434) );
  MUX U1896 ( .IN0(n1502), .IN1(n1503), .SEL(n526), .F(n1499) );
  IV U1897 ( .A(n1504), .Z(n1503) );
  MUX U1898 ( .IN0(n1397), .IN1(n1398), .SEL(iter[3]), .F(n1350) );
  MUX U1899 ( .IN0(n1435), .IN1(n1438), .SEL(n725), .F(n1398) );
  MUX U1900 ( .IN0(n1505), .IN1(n1506), .SEL(iter[1]), .F(n1438) );
  AND U1901 ( .A(n1507), .B(n526), .Z(n1435) );
  MUX U1902 ( .IN0(n1437), .IN1(n1432), .SEL(n725), .F(n1397) );
  MUX U1903 ( .IN0(n1508), .IN1(n1509), .SEL(iter[1]), .F(n1432) );
  MUX U1904 ( .IN0(n1510), .IN1(n1511), .SEL(iter[1]), .F(n1437) );
  IV U1905 ( .A(o[65]), .Z(n1211) );
  XOR U1906 ( .A(n1512), .B(n1513), .Z(n1230) );
  MUX U1907 ( .IN0(n560), .IN1(N36), .SEL(n685), .F(n1513) );
  IV U1908 ( .A(o[31]), .Z(n685) );
  ANDN U1909 ( .A(n1514), .B(iter[5]), .Z(n560) );
  MUX U1910 ( .IN0(n1515), .IN1(n1353), .SEL(iter[4]), .F(n1514) );
  MUX U1911 ( .IN0(n1405), .IN1(n1404), .SEL(n531), .F(n1353) );
  MUX U1912 ( .IN0(n1444), .IN1(n1450), .SEL(iter[2]), .F(n1404) );
  MUX U1913 ( .IN0(n1484), .IN1(n1485), .SEL(iter[1]), .F(n1450) );
  MUX U1914 ( .IN0(o[56]), .IN1(o[55]), .SEL(n528), .F(n1485) );
  MUX U1915 ( .IN0(o[54]), .IN1(o[53]), .SEL(n528), .F(n1484) );
  MUX U1916 ( .IN0(n1473), .IN1(n1483), .SEL(iter[1]), .F(n1444) );
  MUX U1917 ( .IN0(o[52]), .IN1(o[51]), .SEL(n528), .F(n1483) );
  MUX U1918 ( .IN0(o[50]), .IN1(o[49]), .SEL(n528), .F(n1473) );
  MUX U1919 ( .IN0(n1448), .IN1(n1449), .SEL(n725), .F(n1405) );
  MUX U1920 ( .IN0(n1486), .IN1(n1480), .SEL(iter[1]), .F(n1449) );
  MUX U1921 ( .IN0(o[60]), .IN1(o[59]), .SEL(n528), .F(n1480) );
  MUX U1922 ( .IN0(o[58]), .IN1(o[57]), .SEL(n528), .F(n1486) );
  MUX U1923 ( .IN0(n1482), .IN1(n1481), .SEL(n526), .F(n1448) );
  IV U1924 ( .A(iter[1]), .Z(n526) );
  MUX U1925 ( .IN0(o[61]), .IN1(o[62]), .SEL(iter[0]), .F(n1481) );
  AND U1926 ( .A(o[63]), .B(n528), .Z(n1482) );
  MUX U1927 ( .IN0(n1403), .IN1(n1516), .SEL(n531), .F(n1515) );
  IV U1928 ( .A(iter[3]), .Z(n531) );
  MUX U1929 ( .IN0(n1517), .IN1(n1447), .SEL(iter[2]), .F(n1516) );
  MUX U1930 ( .IN0(n1476), .IN1(n1479), .SEL(iter[1]), .F(n1447) );
  MUX U1931 ( .IN0(o[40]), .IN1(o[39]), .SEL(n528), .F(n1479) );
  MUX U1932 ( .IN0(o[38]), .IN1(o[37]), .SEL(n528), .F(n1476) );
  IV U1933 ( .A(n1518), .Z(n1517) );
  MUX U1934 ( .IN0(n1519), .IN1(n1477), .SEL(iter[1]), .F(n1518) );
  MUX U1935 ( .IN0(n917), .IN1(n921), .SEL(iter[0]), .F(n1477) );
  IV U1936 ( .A(o[35]), .Z(n917) );
  MUX U1937 ( .IN0(n913), .IN1(n909), .SEL(n528), .F(n1519) );
  IV U1938 ( .A(o[33]), .Z(n909) );
  IV U1939 ( .A(o[34]), .Z(n913) );
  MUX U1940 ( .IN0(n1446), .IN1(n1445), .SEL(iter[2]), .F(n1403) );
  MUX U1941 ( .IN0(n1471), .IN1(n1472), .SEL(iter[1]), .F(n1445) );
  MUX U1942 ( .IN0(o[48]), .IN1(o[47]), .SEL(n528), .F(n1472) );
  MUX U1943 ( .IN0(o[46]), .IN1(o[45]), .SEL(n528), .F(n1471) );
  MUX U1944 ( .IN0(n1478), .IN1(n1470), .SEL(iter[1]), .F(n1446) );
  MUX U1945 ( .IN0(o[44]), .IN1(o[43]), .SEL(n528), .F(n1470) );
  MUX U1946 ( .IN0(o[42]), .IN1(o[41]), .SEL(n528), .F(n1478) );
  NANDN U1947 ( .B(n1527), .A(o[64]), .Z(n1512) );
  IV U1948 ( .A(n1227), .Z(n1527) );
  AND U1949 ( .A(n1520), .B(n527), .Z(n1227) );
  IV U1950 ( .A(iter[5]), .Z(n527) );
  MUX U1951 ( .IN0(n1356), .IN1(n1521), .SEL(n530), .F(n1520) );
  IV U1952 ( .A(iter[4]), .Z(n530) );
  MUX U1953 ( .IN0(n1522), .IN1(n1410), .SEL(iter[3]), .F(n1521) );
  MUX U1954 ( .IN0(n1457), .IN1(n1523), .SEL(n725), .F(n1410) );
  IV U1955 ( .A(n1459), .Z(n1523) );
  MUX U1956 ( .IN0(n1501), .IN1(n1493), .SEL(iter[1]), .F(n1459) );
  MUX U1957 ( .IN0(n949), .IN1(n945), .SEL(n528), .F(n1493) );
  IV U1958 ( .A(o[42]), .Z(n945) );
  IV U1959 ( .A(o[43]), .Z(n949) );
  MUX U1960 ( .IN0(n941), .IN1(n937), .SEL(n528), .F(n1501) );
  IV U1961 ( .A(o[40]), .Z(n937) );
  IV U1962 ( .A(o[41]), .Z(n941) );
  MUX U1963 ( .IN0(n1495), .IN1(n1496), .SEL(iter[1]), .F(n1457) );
  MUX U1964 ( .IN0(o[46]), .IN1(o[47]), .SEL(iter[0]), .F(n1496) );
  MUX U1965 ( .IN0(o[44]), .IN1(o[45]), .SEL(iter[0]), .F(n1495) );
  MUX U1966 ( .IN0(n1524), .IN1(n1525), .SEL(n725), .F(n1522) );
  IV U1967 ( .A(iter[2]), .Z(n725) );
  MUX U1968 ( .IN0(n1526), .IN1(n1504), .SEL(iter[1]), .F(n1525) );
  MUX U1969 ( .IN0(o[35]), .IN1(o[34]), .SEL(n528), .F(n1504) );
  MUX U1970 ( .IN0(o[33]), .IN1(o[32]), .SEL(n528), .F(n1526) );
  IV U1971 ( .A(n1460), .Z(n1524) );
  MUX U1972 ( .IN0(n1502), .IN1(n1500), .SEL(iter[1]), .F(n1460) );
  MUX U1973 ( .IN0(n933), .IN1(n929), .SEL(n528), .F(n1500) );
  IV U1974 ( .A(o[38]), .Z(n929) );
  IV U1975 ( .A(o[39]), .Z(n933) );
  MUX U1976 ( .IN0(n921), .IN1(n925), .SEL(iter[0]), .F(n1502) );
  IV U1977 ( .A(o[37]), .Z(n925) );
  IV U1978 ( .A(o[36]), .Z(n921) );
  MUX U1979 ( .IN0(n1411), .IN1(n1412), .SEL(iter[3]), .F(n1356) );
  MUX U1980 ( .IN0(n1464), .IN1(n1461), .SEL(iter[2]), .F(n1412) );
  MUX U1981 ( .IN0(n1506), .IN1(n1507), .SEL(iter[1]), .F(n1461) );
  MUX U1982 ( .IN0(o[63]), .IN1(o[62]), .SEL(n528), .F(n1507) );
  MUX U1983 ( .IN0(o[60]), .IN1(o[61]), .SEL(iter[0]), .F(n1506) );
  MUX U1984 ( .IN0(n1511), .IN1(n1505), .SEL(iter[1]), .F(n1464) );
  MUX U1985 ( .IN0(o[59]), .IN1(o[58]), .SEL(n528), .F(n1505) );
  IV U1986 ( .A(iter[0]), .Z(n528) );
  MUX U1987 ( .IN0(o[56]), .IN1(o[57]), .SEL(iter[0]), .F(n1511) );
  MUX U1988 ( .IN0(n1458), .IN1(n1463), .SEL(iter[2]), .F(n1411) );
  MUX U1989 ( .IN0(n1509), .IN1(n1510), .SEL(iter[1]), .F(n1463) );
  MUX U1990 ( .IN0(o[54]), .IN1(o[55]), .SEL(iter[0]), .F(n1510) );
  MUX U1991 ( .IN0(o[52]), .IN1(o[53]), .SEL(iter[0]), .F(n1509) );
  MUX U1992 ( .IN0(n1497), .IN1(n1508), .SEL(iter[1]), .F(n1458) );
  MUX U1993 ( .IN0(o[50]), .IN1(o[51]), .SEL(iter[0]), .F(n1508) );
  MUX U1994 ( .IN0(o[48]), .IN1(o[49]), .SEL(iter[0]), .F(n1497) );
  IV U1995 ( .A(o[94]), .Z(n1299) );
endmodule

