
module matrix_mult_N_M_3_N3_M32 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   \add_24/carry[31] , \add_24/carry[30] , \add_24/carry[29] ,
         \add_24/carry[28] , \add_24/carry[27] , \add_24/carry[26] ,
         \add_24/carry[25] , \add_24/carry[24] , \add_24/carry[23] ,
         \add_24/carry[22] , \add_24/carry[21] , \add_24/carry[20] ,
         \add_24/carry[19] , \add_24/carry[18] , \add_24/carry[17] ,
         \add_24/carry[16] , \add_24/carry[15] , \add_24/carry[14] ,
         \add_24/carry[13] , \add_24/carry[12] , \add_24/carry[11] ,
         \add_24/carry[10] , \add_24/carry[9] , \add_24/carry[8] ,
         \add_24/carry[7] , \add_24/carry[6] , \add_24/carry[5] ,
         \add_24/carry[4] , \add_24/carry[3] , \add_24/carry[2] ,
         \add_24/carry[1] , \mult_23/SUMB[16][1] , \mult_23/SUMB[16][2] ,
         \mult_23/SUMB[16][3] , \mult_23/SUMB[16][4] , \mult_23/SUMB[16][5] ,
         \mult_23/SUMB[16][6] , \mult_23/SUMB[16][7] , \mult_23/SUMB[16][8] ,
         \mult_23/SUMB[16][9] , \mult_23/SUMB[16][10] , \mult_23/SUMB[16][11] ,
         \mult_23/SUMB[16][12] , \mult_23/SUMB[16][13] ,
         \mult_23/SUMB[16][14] , \mult_23/SUMB[16][15] , \mult_23/SUMB[17][1] ,
         \mult_23/SUMB[17][2] , \mult_23/SUMB[17][3] , \mult_23/SUMB[17][4] ,
         \mult_23/SUMB[17][5] , \mult_23/SUMB[17][6] , \mult_23/SUMB[17][7] ,
         \mult_23/SUMB[17][8] , \mult_23/SUMB[17][9] , \mult_23/SUMB[17][10] ,
         \mult_23/SUMB[17][11] , \mult_23/SUMB[17][12] ,
         \mult_23/SUMB[17][13] , \mult_23/SUMB[17][14] , \mult_23/SUMB[18][1] ,
         \mult_23/SUMB[18][2] , \mult_23/SUMB[18][3] , \mult_23/SUMB[18][4] ,
         \mult_23/SUMB[18][5] , \mult_23/SUMB[18][6] , \mult_23/SUMB[18][7] ,
         \mult_23/SUMB[18][8] , \mult_23/SUMB[18][9] , \mult_23/SUMB[18][10] ,
         \mult_23/SUMB[18][11] , \mult_23/SUMB[18][12] ,
         \mult_23/SUMB[18][13] , \mult_23/SUMB[19][1] , \mult_23/SUMB[19][2] ,
         \mult_23/SUMB[19][3] , \mult_23/SUMB[19][4] , \mult_23/SUMB[19][5] ,
         \mult_23/SUMB[19][6] , \mult_23/SUMB[19][7] , \mult_23/SUMB[19][8] ,
         \mult_23/SUMB[19][9] , \mult_23/SUMB[19][10] , \mult_23/SUMB[19][11] ,
         \mult_23/SUMB[19][12] , \mult_23/SUMB[20][1] , \mult_23/SUMB[20][2] ,
         \mult_23/SUMB[20][3] , \mult_23/SUMB[20][4] , \mult_23/SUMB[20][5] ,
         \mult_23/SUMB[20][6] , \mult_23/SUMB[20][7] , \mult_23/SUMB[20][8] ,
         \mult_23/SUMB[20][9] , \mult_23/SUMB[20][10] , \mult_23/SUMB[20][11] ,
         \mult_23/SUMB[21][1] , \mult_23/SUMB[21][2] , \mult_23/SUMB[21][3] ,
         \mult_23/SUMB[21][4] , \mult_23/SUMB[21][5] , \mult_23/SUMB[21][6] ,
         \mult_23/SUMB[21][7] , \mult_23/SUMB[21][8] , \mult_23/SUMB[21][9] ,
         \mult_23/SUMB[21][10] , \mult_23/SUMB[22][1] , \mult_23/SUMB[22][2] ,
         \mult_23/SUMB[22][3] , \mult_23/SUMB[22][4] , \mult_23/SUMB[22][5] ,
         \mult_23/SUMB[22][6] , \mult_23/SUMB[22][7] , \mult_23/SUMB[22][8] ,
         \mult_23/SUMB[22][9] , \mult_23/SUMB[23][1] , \mult_23/SUMB[23][2] ,
         \mult_23/SUMB[23][3] , \mult_23/SUMB[23][4] , \mult_23/SUMB[23][5] ,
         \mult_23/SUMB[23][6] , \mult_23/SUMB[23][7] , \mult_23/SUMB[23][8] ,
         \mult_23/SUMB[24][1] , \mult_23/SUMB[24][2] , \mult_23/SUMB[24][3] ,
         \mult_23/SUMB[24][4] , \mult_23/SUMB[24][5] , \mult_23/SUMB[24][6] ,
         \mult_23/SUMB[24][7] , \mult_23/SUMB[25][1] , \mult_23/SUMB[25][2] ,
         \mult_23/SUMB[25][3] , \mult_23/SUMB[25][4] , \mult_23/SUMB[25][5] ,
         \mult_23/SUMB[25][6] , \mult_23/SUMB[26][1] , \mult_23/SUMB[26][2] ,
         \mult_23/SUMB[26][3] , \mult_23/SUMB[26][4] , \mult_23/SUMB[26][5] ,
         \mult_23/SUMB[27][1] , \mult_23/SUMB[27][2] , \mult_23/SUMB[27][3] ,
         \mult_23/SUMB[27][4] , \mult_23/SUMB[28][1] , \mult_23/SUMB[28][2] ,
         \mult_23/SUMB[28][3] , \mult_23/SUMB[29][1] , \mult_23/SUMB[29][2] ,
         \mult_23/SUMB[30][1] , \mult_23/SUMB[31][0] , \mult_23/CARRYB[16][0] ,
         \mult_23/CARRYB[16][1] , \mult_23/CARRYB[16][2] ,
         \mult_23/CARRYB[16][3] , \mult_23/CARRYB[16][4] ,
         \mult_23/CARRYB[16][5] , \mult_23/CARRYB[16][6] ,
         \mult_23/CARRYB[16][7] , \mult_23/CARRYB[16][8] ,
         \mult_23/CARRYB[16][9] , \mult_23/CARRYB[16][10] ,
         \mult_23/CARRYB[16][11] , \mult_23/CARRYB[16][12] ,
         \mult_23/CARRYB[16][13] , \mult_23/CARRYB[16][14] ,
         \mult_23/CARRYB[17][0] , \mult_23/CARRYB[17][1] ,
         \mult_23/CARRYB[17][2] , \mult_23/CARRYB[17][3] ,
         \mult_23/CARRYB[17][4] , \mult_23/CARRYB[17][5] ,
         \mult_23/CARRYB[17][6] , \mult_23/CARRYB[17][7] ,
         \mult_23/CARRYB[17][8] , \mult_23/CARRYB[17][9] ,
         \mult_23/CARRYB[17][10] , \mult_23/CARRYB[17][11] ,
         \mult_23/CARRYB[17][12] , \mult_23/CARRYB[17][13] ,
         \mult_23/CARRYB[18][0] , \mult_23/CARRYB[18][1] ,
         \mult_23/CARRYB[18][2] , \mult_23/CARRYB[18][3] ,
         \mult_23/CARRYB[18][4] , \mult_23/CARRYB[18][5] ,
         \mult_23/CARRYB[18][6] , \mult_23/CARRYB[18][7] ,
         \mult_23/CARRYB[18][8] , \mult_23/CARRYB[18][9] ,
         \mult_23/CARRYB[18][10] , \mult_23/CARRYB[18][11] ,
         \mult_23/CARRYB[18][12] , \mult_23/CARRYB[19][0] ,
         \mult_23/CARRYB[19][1] , \mult_23/CARRYB[19][2] ,
         \mult_23/CARRYB[19][3] , \mult_23/CARRYB[19][4] ,
         \mult_23/CARRYB[19][5] , \mult_23/CARRYB[19][6] ,
         \mult_23/CARRYB[19][7] , \mult_23/CARRYB[19][8] ,
         \mult_23/CARRYB[19][9] , \mult_23/CARRYB[19][10] ,
         \mult_23/CARRYB[19][11] , \mult_23/CARRYB[20][0] ,
         \mult_23/CARRYB[20][1] , \mult_23/CARRYB[20][2] ,
         \mult_23/CARRYB[20][3] , \mult_23/CARRYB[20][4] ,
         \mult_23/CARRYB[20][5] , \mult_23/CARRYB[20][6] ,
         \mult_23/CARRYB[20][7] , \mult_23/CARRYB[20][8] ,
         \mult_23/CARRYB[20][9] , \mult_23/CARRYB[20][10] ,
         \mult_23/CARRYB[21][0] , \mult_23/CARRYB[21][1] ,
         \mult_23/CARRYB[21][2] , \mult_23/CARRYB[21][3] ,
         \mult_23/CARRYB[21][4] , \mult_23/CARRYB[21][5] ,
         \mult_23/CARRYB[21][6] , \mult_23/CARRYB[21][7] ,
         \mult_23/CARRYB[21][8] , \mult_23/CARRYB[21][9] ,
         \mult_23/CARRYB[22][0] , \mult_23/CARRYB[22][1] ,
         \mult_23/CARRYB[22][2] , \mult_23/CARRYB[22][3] ,
         \mult_23/CARRYB[22][4] , \mult_23/CARRYB[22][5] ,
         \mult_23/CARRYB[22][6] , \mult_23/CARRYB[22][7] ,
         \mult_23/CARRYB[22][8] , \mult_23/CARRYB[23][0] ,
         \mult_23/CARRYB[23][1] , \mult_23/CARRYB[23][2] ,
         \mult_23/CARRYB[23][3] , \mult_23/CARRYB[23][4] ,
         \mult_23/CARRYB[23][5] , \mult_23/CARRYB[23][6] ,
         \mult_23/CARRYB[23][7] , \mult_23/CARRYB[24][0] ,
         \mult_23/CARRYB[24][1] , \mult_23/CARRYB[24][2] ,
         \mult_23/CARRYB[24][3] , \mult_23/CARRYB[24][4] ,
         \mult_23/CARRYB[24][5] , \mult_23/CARRYB[24][6] ,
         \mult_23/CARRYB[25][0] , \mult_23/CARRYB[25][1] ,
         \mult_23/CARRYB[25][2] , \mult_23/CARRYB[25][3] ,
         \mult_23/CARRYB[25][4] , \mult_23/CARRYB[25][5] ,
         \mult_23/CARRYB[26][0] , \mult_23/CARRYB[26][1] ,
         \mult_23/CARRYB[26][2] , \mult_23/CARRYB[26][3] ,
         \mult_23/CARRYB[26][4] , \mult_23/CARRYB[27][0] ,
         \mult_23/CARRYB[27][1] , \mult_23/CARRYB[27][2] ,
         \mult_23/CARRYB[27][3] , \mult_23/CARRYB[28][0] ,
         \mult_23/CARRYB[28][1] , \mult_23/CARRYB[28][2] ,
         \mult_23/CARRYB[29][0] , \mult_23/CARRYB[29][1] ,
         \mult_23/CARRYB[30][0] , \mult_23/SUMB[1][1] , \mult_23/SUMB[1][2] ,
         \mult_23/SUMB[1][3] , \mult_23/SUMB[1][4] , \mult_23/SUMB[1][5] ,
         \mult_23/SUMB[1][6] , \mult_23/SUMB[1][7] , \mult_23/SUMB[1][8] ,
         \mult_23/SUMB[1][9] , \mult_23/SUMB[1][10] , \mult_23/SUMB[1][11] ,
         \mult_23/SUMB[1][12] , \mult_23/SUMB[1][13] , \mult_23/SUMB[1][14] ,
         \mult_23/SUMB[1][15] , \mult_23/SUMB[1][16] , \mult_23/SUMB[1][17] ,
         \mult_23/SUMB[1][18] , \mult_23/SUMB[1][19] , \mult_23/SUMB[1][20] ,
         \mult_23/SUMB[1][21] , \mult_23/SUMB[1][22] , \mult_23/SUMB[1][23] ,
         \mult_23/SUMB[1][24] , \mult_23/SUMB[1][25] , \mult_23/SUMB[1][26] ,
         \mult_23/SUMB[1][27] , \mult_23/SUMB[1][28] , \mult_23/SUMB[1][29] ,
         \mult_23/SUMB[1][30] , \mult_23/SUMB[2][1] , \mult_23/SUMB[2][2] ,
         \mult_23/SUMB[2][3] , \mult_23/SUMB[2][4] , \mult_23/SUMB[2][5] ,
         \mult_23/SUMB[2][6] , \mult_23/SUMB[2][7] , \mult_23/SUMB[2][8] ,
         \mult_23/SUMB[2][9] , \mult_23/SUMB[2][10] , \mult_23/SUMB[2][11] ,
         \mult_23/SUMB[2][12] , \mult_23/SUMB[2][13] , \mult_23/SUMB[2][14] ,
         \mult_23/SUMB[2][15] , \mult_23/SUMB[2][16] , \mult_23/SUMB[2][17] ,
         \mult_23/SUMB[2][18] , \mult_23/SUMB[2][19] , \mult_23/SUMB[2][20] ,
         \mult_23/SUMB[2][21] , \mult_23/SUMB[2][22] , \mult_23/SUMB[2][23] ,
         \mult_23/SUMB[2][24] , \mult_23/SUMB[2][25] , \mult_23/SUMB[2][26] ,
         \mult_23/SUMB[2][27] , \mult_23/SUMB[2][28] , \mult_23/SUMB[2][29] ,
         \mult_23/SUMB[3][1] , \mult_23/SUMB[3][2] , \mult_23/SUMB[3][3] ,
         \mult_23/SUMB[3][4] , \mult_23/SUMB[3][5] , \mult_23/SUMB[3][6] ,
         \mult_23/SUMB[3][7] , \mult_23/SUMB[3][8] , \mult_23/SUMB[3][9] ,
         \mult_23/SUMB[3][10] , \mult_23/SUMB[3][11] , \mult_23/SUMB[3][12] ,
         \mult_23/SUMB[3][13] , \mult_23/SUMB[3][14] , \mult_23/SUMB[3][15] ,
         \mult_23/SUMB[3][16] , \mult_23/SUMB[3][17] , \mult_23/SUMB[3][18] ,
         \mult_23/SUMB[3][19] , \mult_23/SUMB[3][20] , \mult_23/SUMB[3][21] ,
         \mult_23/SUMB[3][22] , \mult_23/SUMB[3][23] , \mult_23/SUMB[3][24] ,
         \mult_23/SUMB[3][25] , \mult_23/SUMB[3][26] , \mult_23/SUMB[3][27] ,
         \mult_23/SUMB[3][28] , \mult_23/SUMB[4][1] , \mult_23/SUMB[4][2] ,
         \mult_23/SUMB[4][3] , \mult_23/SUMB[4][4] , \mult_23/SUMB[4][5] ,
         \mult_23/SUMB[4][6] , \mult_23/SUMB[4][7] , \mult_23/SUMB[4][8] ,
         \mult_23/SUMB[4][9] , \mult_23/SUMB[4][10] , \mult_23/SUMB[4][11] ,
         \mult_23/SUMB[4][12] , \mult_23/SUMB[4][13] , \mult_23/SUMB[4][14] ,
         \mult_23/SUMB[4][15] , \mult_23/SUMB[4][16] , \mult_23/SUMB[4][17] ,
         \mult_23/SUMB[4][18] , \mult_23/SUMB[4][19] , \mult_23/SUMB[4][20] ,
         \mult_23/SUMB[4][21] , \mult_23/SUMB[4][22] , \mult_23/SUMB[4][23] ,
         \mult_23/SUMB[4][24] , \mult_23/SUMB[4][25] , \mult_23/SUMB[4][26] ,
         \mult_23/SUMB[4][27] , \mult_23/SUMB[5][1] , \mult_23/SUMB[5][2] ,
         \mult_23/SUMB[5][3] , \mult_23/SUMB[5][4] , \mult_23/SUMB[5][5] ,
         \mult_23/SUMB[5][6] , \mult_23/SUMB[5][7] , \mult_23/SUMB[5][8] ,
         \mult_23/SUMB[5][9] , \mult_23/SUMB[5][10] , \mult_23/SUMB[5][11] ,
         \mult_23/SUMB[5][12] , \mult_23/SUMB[5][13] , \mult_23/SUMB[5][14] ,
         \mult_23/SUMB[5][15] , \mult_23/SUMB[5][16] , \mult_23/SUMB[5][17] ,
         \mult_23/SUMB[5][18] , \mult_23/SUMB[5][19] , \mult_23/SUMB[5][20] ,
         \mult_23/SUMB[5][21] , \mult_23/SUMB[5][22] , \mult_23/SUMB[5][23] ,
         \mult_23/SUMB[5][24] , \mult_23/SUMB[5][25] , \mult_23/SUMB[5][26] ,
         \mult_23/SUMB[6][1] , \mult_23/SUMB[6][2] , \mult_23/SUMB[6][3] ,
         \mult_23/SUMB[6][4] , \mult_23/SUMB[6][5] , \mult_23/SUMB[6][6] ,
         \mult_23/SUMB[6][7] , \mult_23/SUMB[6][8] , \mult_23/SUMB[6][9] ,
         \mult_23/SUMB[6][10] , \mult_23/SUMB[6][11] , \mult_23/SUMB[6][12] ,
         \mult_23/SUMB[6][13] , \mult_23/SUMB[6][14] , \mult_23/SUMB[6][15] ,
         \mult_23/SUMB[6][16] , \mult_23/SUMB[6][17] , \mult_23/SUMB[6][18] ,
         \mult_23/SUMB[6][19] , \mult_23/SUMB[6][20] , \mult_23/SUMB[6][21] ,
         \mult_23/SUMB[6][22] , \mult_23/SUMB[6][23] , \mult_23/SUMB[6][24] ,
         \mult_23/SUMB[6][25] , \mult_23/SUMB[7][1] , \mult_23/SUMB[7][2] ,
         \mult_23/SUMB[7][3] , \mult_23/SUMB[7][4] , \mult_23/SUMB[7][5] ,
         \mult_23/SUMB[7][6] , \mult_23/SUMB[7][7] , \mult_23/SUMB[7][8] ,
         \mult_23/SUMB[7][9] , \mult_23/SUMB[7][10] , \mult_23/SUMB[7][11] ,
         \mult_23/SUMB[7][12] , \mult_23/SUMB[7][13] , \mult_23/SUMB[7][14] ,
         \mult_23/SUMB[7][15] , \mult_23/SUMB[7][16] , \mult_23/SUMB[7][17] ,
         \mult_23/SUMB[7][18] , \mult_23/SUMB[7][19] , \mult_23/SUMB[7][20] ,
         \mult_23/SUMB[7][21] , \mult_23/SUMB[7][22] , \mult_23/SUMB[7][23] ,
         \mult_23/SUMB[7][24] , \mult_23/SUMB[8][1] , \mult_23/SUMB[8][2] ,
         \mult_23/SUMB[8][3] , \mult_23/SUMB[8][4] , \mult_23/SUMB[8][5] ,
         \mult_23/SUMB[8][6] , \mult_23/SUMB[8][7] , \mult_23/SUMB[8][8] ,
         \mult_23/SUMB[8][9] , \mult_23/SUMB[8][10] , \mult_23/SUMB[8][11] ,
         \mult_23/SUMB[8][12] , \mult_23/SUMB[8][13] , \mult_23/SUMB[8][14] ,
         \mult_23/SUMB[8][15] , \mult_23/SUMB[8][16] , \mult_23/SUMB[8][17] ,
         \mult_23/SUMB[8][18] , \mult_23/SUMB[8][19] , \mult_23/SUMB[8][20] ,
         \mult_23/SUMB[8][21] , \mult_23/SUMB[8][22] , \mult_23/SUMB[8][23] ,
         \mult_23/SUMB[9][1] , \mult_23/SUMB[9][2] , \mult_23/SUMB[9][3] ,
         \mult_23/SUMB[9][4] , \mult_23/SUMB[9][5] , \mult_23/SUMB[9][6] ,
         \mult_23/SUMB[9][7] , \mult_23/SUMB[9][8] , \mult_23/SUMB[9][9] ,
         \mult_23/SUMB[9][10] , \mult_23/SUMB[9][11] , \mult_23/SUMB[9][12] ,
         \mult_23/SUMB[9][13] , \mult_23/SUMB[9][14] , \mult_23/SUMB[9][15] ,
         \mult_23/SUMB[9][16] , \mult_23/SUMB[9][17] , \mult_23/SUMB[9][18] ,
         \mult_23/SUMB[9][19] , \mult_23/SUMB[9][20] , \mult_23/SUMB[9][21] ,
         \mult_23/SUMB[9][22] , \mult_23/SUMB[10][1] , \mult_23/SUMB[10][2] ,
         \mult_23/SUMB[10][3] , \mult_23/SUMB[10][4] , \mult_23/SUMB[10][5] ,
         \mult_23/SUMB[10][6] , \mult_23/SUMB[10][7] , \mult_23/SUMB[10][8] ,
         \mult_23/SUMB[10][9] , \mult_23/SUMB[10][10] , \mult_23/SUMB[10][11] ,
         \mult_23/SUMB[10][12] , \mult_23/SUMB[10][13] ,
         \mult_23/SUMB[10][14] , \mult_23/SUMB[10][15] ,
         \mult_23/SUMB[10][16] , \mult_23/SUMB[10][17] ,
         \mult_23/SUMB[10][18] , \mult_23/SUMB[10][19] ,
         \mult_23/SUMB[10][20] , \mult_23/SUMB[10][21] , \mult_23/SUMB[11][1] ,
         \mult_23/SUMB[11][2] , \mult_23/SUMB[11][3] , \mult_23/SUMB[11][4] ,
         \mult_23/SUMB[11][5] , \mult_23/SUMB[11][6] , \mult_23/SUMB[11][7] ,
         \mult_23/SUMB[11][8] , \mult_23/SUMB[11][9] , \mult_23/SUMB[11][10] ,
         \mult_23/SUMB[11][11] , \mult_23/SUMB[11][12] ,
         \mult_23/SUMB[11][13] , \mult_23/SUMB[11][14] ,
         \mult_23/SUMB[11][15] , \mult_23/SUMB[11][16] ,
         \mult_23/SUMB[11][17] , \mult_23/SUMB[11][18] ,
         \mult_23/SUMB[11][19] , \mult_23/SUMB[11][20] , \mult_23/SUMB[12][1] ,
         \mult_23/SUMB[12][2] , \mult_23/SUMB[12][3] , \mult_23/SUMB[12][4] ,
         \mult_23/SUMB[12][5] , \mult_23/SUMB[12][6] , \mult_23/SUMB[12][7] ,
         \mult_23/SUMB[12][8] , \mult_23/SUMB[12][9] , \mult_23/SUMB[12][10] ,
         \mult_23/SUMB[12][11] , \mult_23/SUMB[12][12] ,
         \mult_23/SUMB[12][13] , \mult_23/SUMB[12][14] ,
         \mult_23/SUMB[12][15] , \mult_23/SUMB[12][16] ,
         \mult_23/SUMB[12][17] , \mult_23/SUMB[12][18] ,
         \mult_23/SUMB[12][19] , \mult_23/SUMB[13][1] , \mult_23/SUMB[13][2] ,
         \mult_23/SUMB[13][3] , \mult_23/SUMB[13][4] , \mult_23/SUMB[13][5] ,
         \mult_23/SUMB[13][6] , \mult_23/SUMB[13][7] , \mult_23/SUMB[13][8] ,
         \mult_23/SUMB[13][9] , \mult_23/SUMB[13][10] , \mult_23/SUMB[13][11] ,
         \mult_23/SUMB[13][12] , \mult_23/SUMB[13][13] ,
         \mult_23/SUMB[13][14] , \mult_23/SUMB[13][15] ,
         \mult_23/SUMB[13][16] , \mult_23/SUMB[13][17] ,
         \mult_23/SUMB[13][18] , \mult_23/SUMB[14][1] , \mult_23/SUMB[14][2] ,
         \mult_23/SUMB[14][3] , \mult_23/SUMB[14][4] , \mult_23/SUMB[14][5] ,
         \mult_23/SUMB[14][6] , \mult_23/SUMB[14][7] , \mult_23/SUMB[14][8] ,
         \mult_23/SUMB[14][9] , \mult_23/SUMB[14][10] , \mult_23/SUMB[14][11] ,
         \mult_23/SUMB[14][12] , \mult_23/SUMB[14][13] ,
         \mult_23/SUMB[14][14] , \mult_23/SUMB[14][15] ,
         \mult_23/SUMB[14][16] , \mult_23/SUMB[14][17] , \mult_23/SUMB[15][1] ,
         \mult_23/SUMB[15][2] , \mult_23/SUMB[15][3] , \mult_23/SUMB[15][4] ,
         \mult_23/SUMB[15][5] , \mult_23/SUMB[15][6] , \mult_23/SUMB[15][7] ,
         \mult_23/SUMB[15][8] , \mult_23/SUMB[15][9] , \mult_23/SUMB[15][10] ,
         \mult_23/SUMB[15][11] , \mult_23/SUMB[15][12] ,
         \mult_23/SUMB[15][13] , \mult_23/SUMB[15][14] ,
         \mult_23/SUMB[15][15] , \mult_23/SUMB[15][16] ,
         \mult_23/CARRYB[1][0] , \mult_23/CARRYB[1][1] ,
         \mult_23/CARRYB[1][2] , \mult_23/CARRYB[1][3] ,
         \mult_23/CARRYB[1][4] , \mult_23/CARRYB[1][5] ,
         \mult_23/CARRYB[1][6] , \mult_23/CARRYB[1][7] ,
         \mult_23/CARRYB[1][8] , \mult_23/CARRYB[1][9] ,
         \mult_23/CARRYB[1][10] , \mult_23/CARRYB[1][11] ,
         \mult_23/CARRYB[1][12] , \mult_23/CARRYB[1][13] ,
         \mult_23/CARRYB[1][14] , \mult_23/CARRYB[1][15] ,
         \mult_23/CARRYB[1][16] , \mult_23/CARRYB[1][17] ,
         \mult_23/CARRYB[1][18] , \mult_23/CARRYB[1][19] ,
         \mult_23/CARRYB[1][20] , \mult_23/CARRYB[1][21] ,
         \mult_23/CARRYB[1][22] , \mult_23/CARRYB[1][23] ,
         \mult_23/CARRYB[1][24] , \mult_23/CARRYB[1][25] ,
         \mult_23/CARRYB[1][26] , \mult_23/CARRYB[1][27] ,
         \mult_23/CARRYB[1][28] , \mult_23/CARRYB[1][29] ,
         \mult_23/CARRYB[2][0] , \mult_23/CARRYB[2][1] ,
         \mult_23/CARRYB[2][2] , \mult_23/CARRYB[2][3] ,
         \mult_23/CARRYB[2][4] , \mult_23/CARRYB[2][5] ,
         \mult_23/CARRYB[2][6] , \mult_23/CARRYB[2][7] ,
         \mult_23/CARRYB[2][8] , \mult_23/CARRYB[2][9] ,
         \mult_23/CARRYB[2][10] , \mult_23/CARRYB[2][11] ,
         \mult_23/CARRYB[2][12] , \mult_23/CARRYB[2][13] ,
         \mult_23/CARRYB[2][14] , \mult_23/CARRYB[2][15] ,
         \mult_23/CARRYB[2][16] , \mult_23/CARRYB[2][17] ,
         \mult_23/CARRYB[2][18] , \mult_23/CARRYB[2][19] ,
         \mult_23/CARRYB[2][20] , \mult_23/CARRYB[2][21] ,
         \mult_23/CARRYB[2][22] , \mult_23/CARRYB[2][23] ,
         \mult_23/CARRYB[2][24] , \mult_23/CARRYB[2][25] ,
         \mult_23/CARRYB[2][26] , \mult_23/CARRYB[2][27] ,
         \mult_23/CARRYB[2][28] , \mult_23/CARRYB[3][0] ,
         \mult_23/CARRYB[3][1] , \mult_23/CARRYB[3][2] ,
         \mult_23/CARRYB[3][3] , \mult_23/CARRYB[3][4] ,
         \mult_23/CARRYB[3][5] , \mult_23/CARRYB[3][6] ,
         \mult_23/CARRYB[3][7] , \mult_23/CARRYB[3][8] ,
         \mult_23/CARRYB[3][9] , \mult_23/CARRYB[3][10] ,
         \mult_23/CARRYB[3][11] , \mult_23/CARRYB[3][12] ,
         \mult_23/CARRYB[3][13] , \mult_23/CARRYB[3][14] ,
         \mult_23/CARRYB[3][15] , \mult_23/CARRYB[3][16] ,
         \mult_23/CARRYB[3][17] , \mult_23/CARRYB[3][18] ,
         \mult_23/CARRYB[3][19] , \mult_23/CARRYB[3][20] ,
         \mult_23/CARRYB[3][21] , \mult_23/CARRYB[3][22] ,
         \mult_23/CARRYB[3][23] , \mult_23/CARRYB[3][24] ,
         \mult_23/CARRYB[3][25] , \mult_23/CARRYB[3][26] ,
         \mult_23/CARRYB[3][27] , \mult_23/CARRYB[4][0] ,
         \mult_23/CARRYB[4][1] , \mult_23/CARRYB[4][2] ,
         \mult_23/CARRYB[4][3] , \mult_23/CARRYB[4][4] ,
         \mult_23/CARRYB[4][5] , \mult_23/CARRYB[4][6] ,
         \mult_23/CARRYB[4][7] , \mult_23/CARRYB[4][8] ,
         \mult_23/CARRYB[4][9] , \mult_23/CARRYB[4][10] ,
         \mult_23/CARRYB[4][11] , \mult_23/CARRYB[4][12] ,
         \mult_23/CARRYB[4][13] , \mult_23/CARRYB[4][14] ,
         \mult_23/CARRYB[4][15] , \mult_23/CARRYB[4][16] ,
         \mult_23/CARRYB[4][17] , \mult_23/CARRYB[4][18] ,
         \mult_23/CARRYB[4][19] , \mult_23/CARRYB[4][20] ,
         \mult_23/CARRYB[4][21] , \mult_23/CARRYB[4][22] ,
         \mult_23/CARRYB[4][23] , \mult_23/CARRYB[4][24] ,
         \mult_23/CARRYB[4][25] , \mult_23/CARRYB[4][26] ,
         \mult_23/CARRYB[5][0] , \mult_23/CARRYB[5][1] ,
         \mult_23/CARRYB[5][2] , \mult_23/CARRYB[5][3] ,
         \mult_23/CARRYB[5][4] , \mult_23/CARRYB[5][5] ,
         \mult_23/CARRYB[5][6] , \mult_23/CARRYB[5][7] ,
         \mult_23/CARRYB[5][8] , \mult_23/CARRYB[5][9] ,
         \mult_23/CARRYB[5][10] , \mult_23/CARRYB[5][11] ,
         \mult_23/CARRYB[5][12] , \mult_23/CARRYB[5][13] ,
         \mult_23/CARRYB[5][14] , \mult_23/CARRYB[5][15] ,
         \mult_23/CARRYB[5][16] , \mult_23/CARRYB[5][17] ,
         \mult_23/CARRYB[5][18] , \mult_23/CARRYB[5][19] ,
         \mult_23/CARRYB[5][20] , \mult_23/CARRYB[5][21] ,
         \mult_23/CARRYB[5][22] , \mult_23/CARRYB[5][23] ,
         \mult_23/CARRYB[5][24] , \mult_23/CARRYB[5][25] ,
         \mult_23/CARRYB[6][0] , \mult_23/CARRYB[6][1] ,
         \mult_23/CARRYB[6][2] , \mult_23/CARRYB[6][3] ,
         \mult_23/CARRYB[6][4] , \mult_23/CARRYB[6][5] ,
         \mult_23/CARRYB[6][6] , \mult_23/CARRYB[6][7] ,
         \mult_23/CARRYB[6][8] , \mult_23/CARRYB[6][9] ,
         \mult_23/CARRYB[6][10] , \mult_23/CARRYB[6][11] ,
         \mult_23/CARRYB[6][12] , \mult_23/CARRYB[6][13] ,
         \mult_23/CARRYB[6][14] , \mult_23/CARRYB[6][15] ,
         \mult_23/CARRYB[6][16] , \mult_23/CARRYB[6][17] ,
         \mult_23/CARRYB[6][18] , \mult_23/CARRYB[6][19] ,
         \mult_23/CARRYB[6][20] , \mult_23/CARRYB[6][21] ,
         \mult_23/CARRYB[6][22] , \mult_23/CARRYB[6][23] ,
         \mult_23/CARRYB[6][24] , \mult_23/CARRYB[7][0] ,
         \mult_23/CARRYB[7][1] , \mult_23/CARRYB[7][2] ,
         \mult_23/CARRYB[7][3] , \mult_23/CARRYB[7][4] ,
         \mult_23/CARRYB[7][5] , \mult_23/CARRYB[7][6] ,
         \mult_23/CARRYB[7][7] , \mult_23/CARRYB[7][8] ,
         \mult_23/CARRYB[7][9] , \mult_23/CARRYB[7][10] ,
         \mult_23/CARRYB[7][11] , \mult_23/CARRYB[7][12] ,
         \mult_23/CARRYB[7][13] , \mult_23/CARRYB[7][14] ,
         \mult_23/CARRYB[7][15] , \mult_23/CARRYB[7][16] ,
         \mult_23/CARRYB[7][17] , \mult_23/CARRYB[7][18] ,
         \mult_23/CARRYB[7][19] , \mult_23/CARRYB[7][20] ,
         \mult_23/CARRYB[7][21] , \mult_23/CARRYB[7][22] ,
         \mult_23/CARRYB[7][23] , \mult_23/CARRYB[8][0] ,
         \mult_23/CARRYB[8][1] , \mult_23/CARRYB[8][2] ,
         \mult_23/CARRYB[8][3] , \mult_23/CARRYB[8][4] ,
         \mult_23/CARRYB[8][5] , \mult_23/CARRYB[8][6] ,
         \mult_23/CARRYB[8][7] , \mult_23/CARRYB[8][8] ,
         \mult_23/CARRYB[8][9] , \mult_23/CARRYB[8][10] ,
         \mult_23/CARRYB[8][11] , \mult_23/CARRYB[8][12] ,
         \mult_23/CARRYB[8][13] , \mult_23/CARRYB[8][14] ,
         \mult_23/CARRYB[8][15] , \mult_23/CARRYB[8][16] ,
         \mult_23/CARRYB[8][17] , \mult_23/CARRYB[8][18] ,
         \mult_23/CARRYB[8][19] , \mult_23/CARRYB[8][20] ,
         \mult_23/CARRYB[8][21] , \mult_23/CARRYB[8][22] ,
         \mult_23/CARRYB[9][0] , \mult_23/CARRYB[9][1] ,
         \mult_23/CARRYB[9][2] , \mult_23/CARRYB[9][3] ,
         \mult_23/CARRYB[9][4] , \mult_23/CARRYB[9][5] ,
         \mult_23/CARRYB[9][6] , \mult_23/CARRYB[9][7] ,
         \mult_23/CARRYB[9][8] , \mult_23/CARRYB[9][9] ,
         \mult_23/CARRYB[9][10] , \mult_23/CARRYB[9][11] ,
         \mult_23/CARRYB[9][12] , \mult_23/CARRYB[9][13] ,
         \mult_23/CARRYB[9][14] , \mult_23/CARRYB[9][15] ,
         \mult_23/CARRYB[9][16] , \mult_23/CARRYB[9][17] ,
         \mult_23/CARRYB[9][18] , \mult_23/CARRYB[9][19] ,
         \mult_23/CARRYB[9][20] , \mult_23/CARRYB[9][21] ,
         \mult_23/CARRYB[10][0] , \mult_23/CARRYB[10][1] ,
         \mult_23/CARRYB[10][2] , \mult_23/CARRYB[10][3] ,
         \mult_23/CARRYB[10][4] , \mult_23/CARRYB[10][5] ,
         \mult_23/CARRYB[10][6] , \mult_23/CARRYB[10][7] ,
         \mult_23/CARRYB[10][8] , \mult_23/CARRYB[10][9] ,
         \mult_23/CARRYB[10][10] , \mult_23/CARRYB[10][11] ,
         \mult_23/CARRYB[10][12] , \mult_23/CARRYB[10][13] ,
         \mult_23/CARRYB[10][14] , \mult_23/CARRYB[10][15] ,
         \mult_23/CARRYB[10][16] , \mult_23/CARRYB[10][17] ,
         \mult_23/CARRYB[10][18] , \mult_23/CARRYB[10][19] ,
         \mult_23/CARRYB[10][20] , \mult_23/CARRYB[11][0] ,
         \mult_23/CARRYB[11][1] , \mult_23/CARRYB[11][2] ,
         \mult_23/CARRYB[11][3] , \mult_23/CARRYB[11][4] ,
         \mult_23/CARRYB[11][5] , \mult_23/CARRYB[11][6] ,
         \mult_23/CARRYB[11][7] , \mult_23/CARRYB[11][8] ,
         \mult_23/CARRYB[11][9] , \mult_23/CARRYB[11][10] ,
         \mult_23/CARRYB[11][11] , \mult_23/CARRYB[11][12] ,
         \mult_23/CARRYB[11][13] , \mult_23/CARRYB[11][14] ,
         \mult_23/CARRYB[11][15] , \mult_23/CARRYB[11][16] ,
         \mult_23/CARRYB[11][17] , \mult_23/CARRYB[11][18] ,
         \mult_23/CARRYB[11][19] , \mult_23/CARRYB[12][0] ,
         \mult_23/CARRYB[12][1] , \mult_23/CARRYB[12][2] ,
         \mult_23/CARRYB[12][3] , \mult_23/CARRYB[12][4] ,
         \mult_23/CARRYB[12][5] , \mult_23/CARRYB[12][6] ,
         \mult_23/CARRYB[12][7] , \mult_23/CARRYB[12][8] ,
         \mult_23/CARRYB[12][9] , \mult_23/CARRYB[12][10] ,
         \mult_23/CARRYB[12][11] , \mult_23/CARRYB[12][12] ,
         \mult_23/CARRYB[12][13] , \mult_23/CARRYB[12][14] ,
         \mult_23/CARRYB[12][15] , \mult_23/CARRYB[12][16] ,
         \mult_23/CARRYB[12][17] , \mult_23/CARRYB[12][18] ,
         \mult_23/CARRYB[13][0] , \mult_23/CARRYB[13][1] ,
         \mult_23/CARRYB[13][2] , \mult_23/CARRYB[13][3] ,
         \mult_23/CARRYB[13][4] , \mult_23/CARRYB[13][5] ,
         \mult_23/CARRYB[13][6] , \mult_23/CARRYB[13][7] ,
         \mult_23/CARRYB[13][8] , \mult_23/CARRYB[13][9] ,
         \mult_23/CARRYB[13][10] , \mult_23/CARRYB[13][11] ,
         \mult_23/CARRYB[13][12] , \mult_23/CARRYB[13][13] ,
         \mult_23/CARRYB[13][14] , \mult_23/CARRYB[13][15] ,
         \mult_23/CARRYB[13][16] , \mult_23/CARRYB[13][17] ,
         \mult_23/CARRYB[14][0] , \mult_23/CARRYB[14][1] ,
         \mult_23/CARRYB[14][2] , \mult_23/CARRYB[14][3] ,
         \mult_23/CARRYB[14][4] , \mult_23/CARRYB[14][5] ,
         \mult_23/CARRYB[14][6] , \mult_23/CARRYB[14][7] ,
         \mult_23/CARRYB[14][8] , \mult_23/CARRYB[14][9] ,
         \mult_23/CARRYB[14][10] , \mult_23/CARRYB[14][11] ,
         \mult_23/CARRYB[14][12] , \mult_23/CARRYB[14][13] ,
         \mult_23/CARRYB[14][14] , \mult_23/CARRYB[14][15] ,
         \mult_23/CARRYB[14][16] , \mult_23/CARRYB[15][0] ,
         \mult_23/CARRYB[15][1] , \mult_23/CARRYB[15][2] ,
         \mult_23/CARRYB[15][3] , \mult_23/CARRYB[15][4] ,
         \mult_23/CARRYB[15][5] , \mult_23/CARRYB[15][6] ,
         \mult_23/CARRYB[15][7] , \mult_23/CARRYB[15][8] ,
         \mult_23/CARRYB[15][9] , \mult_23/CARRYB[15][10] ,
         \mult_23/CARRYB[15][11] , \mult_23/CARRYB[15][12] ,
         \mult_23/CARRYB[15][13] , \mult_23/CARRYB[15][14] ,
         \mult_23/CARRYB[15][15] , \mult_23/ab[0][1] , \mult_23/ab[0][2] ,
         \mult_23/ab[0][3] , \mult_23/ab[0][4] , \mult_23/ab[0][5] ,
         \mult_23/ab[0][6] , \mult_23/ab[0][7] , \mult_23/ab[0][8] ,
         \mult_23/ab[0][9] , \mult_23/ab[0][10] , \mult_23/ab[0][11] ,
         \mult_23/ab[0][12] , \mult_23/ab[0][13] , \mult_23/ab[0][14] ,
         \mult_23/ab[0][15] , \mult_23/ab[0][16] , \mult_23/ab[0][17] ,
         \mult_23/ab[0][18] , \mult_23/ab[0][19] , \mult_23/ab[0][20] ,
         \mult_23/ab[0][21] , \mult_23/ab[0][22] , \mult_23/ab[0][23] ,
         \mult_23/ab[0][24] , \mult_23/ab[0][25] , \mult_23/ab[0][26] ,
         \mult_23/ab[0][27] , \mult_23/ab[0][28] , \mult_23/ab[0][29] ,
         \mult_23/ab[0][30] , \mult_23/ab[0][31] , \mult_23/ab[1][0] ,
         \mult_23/ab[1][1] , \mult_23/ab[1][2] , \mult_23/ab[1][3] ,
         \mult_23/ab[1][4] , \mult_23/ab[1][5] , \mult_23/ab[1][6] ,
         \mult_23/ab[1][7] , \mult_23/ab[1][8] , \mult_23/ab[1][9] ,
         \mult_23/ab[1][10] , \mult_23/ab[1][11] , \mult_23/ab[1][12] ,
         \mult_23/ab[1][13] , \mult_23/ab[1][14] , \mult_23/ab[1][15] ,
         \mult_23/ab[1][16] , \mult_23/ab[1][17] , \mult_23/ab[1][18] ,
         \mult_23/ab[1][19] , \mult_23/ab[1][20] , \mult_23/ab[1][21] ,
         \mult_23/ab[1][22] , \mult_23/ab[1][23] , \mult_23/ab[1][24] ,
         \mult_23/ab[1][25] , \mult_23/ab[1][26] , \mult_23/ab[1][27] ,
         \mult_23/ab[1][28] , \mult_23/ab[1][29] , \mult_23/ab[1][30] ,
         \mult_23/ab[2][0] , \mult_23/ab[2][1] , \mult_23/ab[2][2] ,
         \mult_23/ab[2][3] , \mult_23/ab[2][4] , \mult_23/ab[2][5] ,
         \mult_23/ab[2][6] , \mult_23/ab[2][7] , \mult_23/ab[2][8] ,
         \mult_23/ab[2][9] , \mult_23/ab[2][10] , \mult_23/ab[2][11] ,
         \mult_23/ab[2][12] , \mult_23/ab[2][13] , \mult_23/ab[2][14] ,
         \mult_23/ab[2][15] , \mult_23/ab[2][16] , \mult_23/ab[2][17] ,
         \mult_23/ab[2][18] , \mult_23/ab[2][19] , \mult_23/ab[2][20] ,
         \mult_23/ab[2][21] , \mult_23/ab[2][22] , \mult_23/ab[2][23] ,
         \mult_23/ab[2][24] , \mult_23/ab[2][25] , \mult_23/ab[2][26] ,
         \mult_23/ab[2][27] , \mult_23/ab[2][28] , \mult_23/ab[2][29] ,
         \mult_23/ab[3][0] , \mult_23/ab[3][1] , \mult_23/ab[3][2] ,
         \mult_23/ab[3][3] , \mult_23/ab[3][4] , \mult_23/ab[3][5] ,
         \mult_23/ab[3][6] , \mult_23/ab[3][7] , \mult_23/ab[3][8] ,
         \mult_23/ab[3][9] , \mult_23/ab[3][10] , \mult_23/ab[3][11] ,
         \mult_23/ab[3][12] , \mult_23/ab[3][13] , \mult_23/ab[3][14] ,
         \mult_23/ab[3][15] , \mult_23/ab[3][16] , \mult_23/ab[3][17] ,
         \mult_23/ab[3][18] , \mult_23/ab[3][19] , \mult_23/ab[3][20] ,
         \mult_23/ab[3][21] , \mult_23/ab[3][22] , \mult_23/ab[3][23] ,
         \mult_23/ab[3][24] , \mult_23/ab[3][25] , \mult_23/ab[3][26] ,
         \mult_23/ab[3][27] , \mult_23/ab[3][28] , \mult_23/ab[4][0] ,
         \mult_23/ab[4][1] , \mult_23/ab[4][2] , \mult_23/ab[4][3] ,
         \mult_23/ab[4][4] , \mult_23/ab[4][5] , \mult_23/ab[4][6] ,
         \mult_23/ab[4][7] , \mult_23/ab[4][8] , \mult_23/ab[4][9] ,
         \mult_23/ab[4][10] , \mult_23/ab[4][11] , \mult_23/ab[4][12] ,
         \mult_23/ab[4][13] , \mult_23/ab[4][14] , \mult_23/ab[4][15] ,
         \mult_23/ab[4][16] , \mult_23/ab[4][17] , \mult_23/ab[4][18] ,
         \mult_23/ab[4][19] , \mult_23/ab[4][20] , \mult_23/ab[4][21] ,
         \mult_23/ab[4][22] , \mult_23/ab[4][23] , \mult_23/ab[4][24] ,
         \mult_23/ab[4][25] , \mult_23/ab[4][26] , \mult_23/ab[4][27] ,
         \mult_23/ab[5][0] , \mult_23/ab[5][1] , \mult_23/ab[5][2] ,
         \mult_23/ab[5][3] , \mult_23/ab[5][4] , \mult_23/ab[5][5] ,
         \mult_23/ab[5][6] , \mult_23/ab[5][7] , \mult_23/ab[5][8] ,
         \mult_23/ab[5][9] , \mult_23/ab[5][10] , \mult_23/ab[5][11] ,
         \mult_23/ab[5][12] , \mult_23/ab[5][13] , \mult_23/ab[5][14] ,
         \mult_23/ab[5][15] , \mult_23/ab[5][16] , \mult_23/ab[5][17] ,
         \mult_23/ab[5][18] , \mult_23/ab[5][19] , \mult_23/ab[5][20] ,
         \mult_23/ab[5][21] , \mult_23/ab[5][22] , \mult_23/ab[5][23] ,
         \mult_23/ab[5][24] , \mult_23/ab[5][25] , \mult_23/ab[5][26] ,
         \mult_23/ab[6][0] , \mult_23/ab[6][1] , \mult_23/ab[6][2] ,
         \mult_23/ab[6][3] , \mult_23/ab[6][4] , \mult_23/ab[6][5] ,
         \mult_23/ab[6][6] , \mult_23/ab[6][7] , \mult_23/ab[6][8] ,
         \mult_23/ab[6][9] , \mult_23/ab[6][10] , \mult_23/ab[6][11] ,
         \mult_23/ab[6][12] , \mult_23/ab[6][13] , \mult_23/ab[6][14] ,
         \mult_23/ab[6][15] , \mult_23/ab[6][16] , \mult_23/ab[6][17] ,
         \mult_23/ab[6][18] , \mult_23/ab[6][19] , \mult_23/ab[6][20] ,
         \mult_23/ab[6][21] , \mult_23/ab[6][22] , \mult_23/ab[6][23] ,
         \mult_23/ab[6][24] , \mult_23/ab[6][25] , \mult_23/ab[7][0] ,
         \mult_23/ab[7][1] , \mult_23/ab[7][2] , \mult_23/ab[7][3] ,
         \mult_23/ab[7][4] , \mult_23/ab[7][5] , \mult_23/ab[7][6] ,
         \mult_23/ab[7][7] , \mult_23/ab[7][8] , \mult_23/ab[7][9] ,
         \mult_23/ab[7][10] , \mult_23/ab[7][11] , \mult_23/ab[7][12] ,
         \mult_23/ab[7][13] , \mult_23/ab[7][14] , \mult_23/ab[7][15] ,
         \mult_23/ab[7][16] , \mult_23/ab[7][17] , \mult_23/ab[7][18] ,
         \mult_23/ab[7][19] , \mult_23/ab[7][20] , \mult_23/ab[7][21] ,
         \mult_23/ab[7][22] , \mult_23/ab[7][23] , \mult_23/ab[7][24] ,
         \mult_23/ab[8][0] , \mult_23/ab[8][1] , \mult_23/ab[8][2] ,
         \mult_23/ab[8][3] , \mult_23/ab[8][4] , \mult_23/ab[8][5] ,
         \mult_23/ab[8][6] , \mult_23/ab[8][7] , \mult_23/ab[8][8] ,
         \mult_23/ab[8][9] , \mult_23/ab[8][10] , \mult_23/ab[8][11] ,
         \mult_23/ab[8][12] , \mult_23/ab[8][13] , \mult_23/ab[8][14] ,
         \mult_23/ab[8][15] , \mult_23/ab[8][16] , \mult_23/ab[8][17] ,
         \mult_23/ab[8][18] , \mult_23/ab[8][19] , \mult_23/ab[8][20] ,
         \mult_23/ab[8][21] , \mult_23/ab[8][22] , \mult_23/ab[8][23] ,
         \mult_23/ab[9][0] , \mult_23/ab[9][1] , \mult_23/ab[9][2] ,
         \mult_23/ab[9][3] , \mult_23/ab[9][4] , \mult_23/ab[9][5] ,
         \mult_23/ab[9][6] , \mult_23/ab[9][7] , \mult_23/ab[9][8] ,
         \mult_23/ab[9][9] , \mult_23/ab[9][10] , \mult_23/ab[9][11] ,
         \mult_23/ab[9][12] , \mult_23/ab[9][13] , \mult_23/ab[9][14] ,
         \mult_23/ab[9][15] , \mult_23/ab[9][16] , \mult_23/ab[9][17] ,
         \mult_23/ab[9][18] , \mult_23/ab[9][19] , \mult_23/ab[9][20] ,
         \mult_23/ab[9][21] , \mult_23/ab[9][22] , \mult_23/ab[10][0] ,
         \mult_23/ab[10][1] , \mult_23/ab[10][2] , \mult_23/ab[10][3] ,
         \mult_23/ab[10][4] , \mult_23/ab[10][5] , \mult_23/ab[10][6] ,
         \mult_23/ab[10][7] , \mult_23/ab[10][8] , \mult_23/ab[10][9] ,
         \mult_23/ab[10][10] , \mult_23/ab[10][11] , \mult_23/ab[10][12] ,
         \mult_23/ab[10][13] , \mult_23/ab[10][14] , \mult_23/ab[10][15] ,
         \mult_23/ab[10][16] , \mult_23/ab[10][17] , \mult_23/ab[10][18] ,
         \mult_23/ab[10][19] , \mult_23/ab[10][20] , \mult_23/ab[10][21] ,
         \mult_23/ab[11][0] , \mult_23/ab[11][1] , \mult_23/ab[11][2] ,
         \mult_23/ab[11][3] , \mult_23/ab[11][4] , \mult_23/ab[11][5] ,
         \mult_23/ab[11][6] , \mult_23/ab[11][7] , \mult_23/ab[11][8] ,
         \mult_23/ab[11][9] , \mult_23/ab[11][10] , \mult_23/ab[11][11] ,
         \mult_23/ab[11][12] , \mult_23/ab[11][13] , \mult_23/ab[11][14] ,
         \mult_23/ab[11][15] , \mult_23/ab[11][16] , \mult_23/ab[11][17] ,
         \mult_23/ab[11][18] , \mult_23/ab[11][19] , \mult_23/ab[11][20] ,
         \mult_23/ab[12][0] , \mult_23/ab[12][1] , \mult_23/ab[12][2] ,
         \mult_23/ab[12][3] , \mult_23/ab[12][4] , \mult_23/ab[12][5] ,
         \mult_23/ab[12][6] , \mult_23/ab[12][7] , \mult_23/ab[12][8] ,
         \mult_23/ab[12][9] , \mult_23/ab[12][10] , \mult_23/ab[12][11] ,
         \mult_23/ab[12][12] , \mult_23/ab[12][13] , \mult_23/ab[12][14] ,
         \mult_23/ab[12][15] , \mult_23/ab[12][16] , \mult_23/ab[12][17] ,
         \mult_23/ab[12][18] , \mult_23/ab[12][19] , \mult_23/ab[13][0] ,
         \mult_23/ab[13][1] , \mult_23/ab[13][2] , \mult_23/ab[13][3] ,
         \mult_23/ab[13][4] , \mult_23/ab[13][5] , \mult_23/ab[13][6] ,
         \mult_23/ab[13][7] , \mult_23/ab[13][8] , \mult_23/ab[13][9] ,
         \mult_23/ab[13][10] , \mult_23/ab[13][11] , \mult_23/ab[13][12] ,
         \mult_23/ab[13][13] , \mult_23/ab[13][14] , \mult_23/ab[13][15] ,
         \mult_23/ab[13][16] , \mult_23/ab[13][17] , \mult_23/ab[13][18] ,
         \mult_23/ab[14][0] , \mult_23/ab[14][1] , \mult_23/ab[14][2] ,
         \mult_23/ab[14][3] , \mult_23/ab[14][4] , \mult_23/ab[14][5] ,
         \mult_23/ab[14][6] , \mult_23/ab[14][7] , \mult_23/ab[14][8] ,
         \mult_23/ab[14][9] , \mult_23/ab[14][10] , \mult_23/ab[14][11] ,
         \mult_23/ab[14][12] , \mult_23/ab[14][13] , \mult_23/ab[14][14] ,
         \mult_23/ab[14][15] , \mult_23/ab[14][16] , \mult_23/ab[14][17] ,
         \mult_23/ab[15][0] , \mult_23/ab[15][1] , \mult_23/ab[15][2] ,
         \mult_23/ab[15][3] , \mult_23/ab[15][4] , \mult_23/ab[15][5] ,
         \mult_23/ab[15][6] , \mult_23/ab[15][7] , \mult_23/ab[15][8] ,
         \mult_23/ab[15][9] , \mult_23/ab[15][10] , \mult_23/ab[15][11] ,
         \mult_23/ab[15][12] , \mult_23/ab[15][13] , \mult_23/ab[15][14] ,
         \mult_23/ab[15][15] , \mult_23/ab[15][16] , \mult_23/ab[16][0] ,
         \mult_23/ab[16][1] , \mult_23/ab[16][2] , \mult_23/ab[16][3] ,
         \mult_23/ab[16][4] , \mult_23/ab[16][5] , \mult_23/ab[16][6] ,
         \mult_23/ab[16][7] , \mult_23/ab[16][8] , \mult_23/ab[16][9] ,
         \mult_23/ab[16][10] , \mult_23/ab[16][11] , \mult_23/ab[16][12] ,
         \mult_23/ab[16][13] , \mult_23/ab[16][14] , \mult_23/ab[16][15] ,
         \mult_23/ab[17][0] , \mult_23/ab[17][1] , \mult_23/ab[17][2] ,
         \mult_23/ab[17][3] , \mult_23/ab[17][4] , \mult_23/ab[17][5] ,
         \mult_23/ab[17][6] , \mult_23/ab[17][7] , \mult_23/ab[17][8] ,
         \mult_23/ab[17][9] , \mult_23/ab[17][10] , \mult_23/ab[17][11] ,
         \mult_23/ab[17][12] , \mult_23/ab[17][13] , \mult_23/ab[17][14] ,
         \mult_23/ab[18][0] , \mult_23/ab[18][1] , \mult_23/ab[18][2] ,
         \mult_23/ab[18][3] , \mult_23/ab[18][4] , \mult_23/ab[18][5] ,
         \mult_23/ab[18][6] , \mult_23/ab[18][7] , \mult_23/ab[18][8] ,
         \mult_23/ab[18][9] , \mult_23/ab[18][10] , \mult_23/ab[18][11] ,
         \mult_23/ab[18][12] , \mult_23/ab[18][13] , \mult_23/ab[19][0] ,
         \mult_23/ab[19][1] , \mult_23/ab[19][2] , \mult_23/ab[19][3] ,
         \mult_23/ab[19][4] , \mult_23/ab[19][5] , \mult_23/ab[19][6] ,
         \mult_23/ab[19][7] , \mult_23/ab[19][8] , \mult_23/ab[19][9] ,
         \mult_23/ab[19][10] , \mult_23/ab[19][11] , \mult_23/ab[19][12] ,
         \mult_23/ab[20][0] , \mult_23/ab[20][1] , \mult_23/ab[20][2] ,
         \mult_23/ab[20][3] , \mult_23/ab[20][4] , \mult_23/ab[20][5] ,
         \mult_23/ab[20][6] , \mult_23/ab[20][7] , \mult_23/ab[20][8] ,
         \mult_23/ab[20][9] , \mult_23/ab[20][10] , \mult_23/ab[20][11] ,
         \mult_23/ab[21][0] , \mult_23/ab[21][1] , \mult_23/ab[21][2] ,
         \mult_23/ab[21][3] , \mult_23/ab[21][4] , \mult_23/ab[21][5] ,
         \mult_23/ab[21][6] , \mult_23/ab[21][7] , \mult_23/ab[21][8] ,
         \mult_23/ab[21][9] , \mult_23/ab[21][10] , \mult_23/ab[22][0] ,
         \mult_23/ab[22][1] , \mult_23/ab[22][2] , \mult_23/ab[22][3] ,
         \mult_23/ab[22][4] , \mult_23/ab[22][5] , \mult_23/ab[22][6] ,
         \mult_23/ab[22][7] , \mult_23/ab[22][8] , \mult_23/ab[22][9] ,
         \mult_23/ab[23][0] , \mult_23/ab[23][1] , \mult_23/ab[23][2] ,
         \mult_23/ab[23][3] , \mult_23/ab[23][4] , \mult_23/ab[23][5] ,
         \mult_23/ab[23][6] , \mult_23/ab[23][7] , \mult_23/ab[23][8] ,
         \mult_23/ab[24][0] , \mult_23/ab[24][1] , \mult_23/ab[24][2] ,
         \mult_23/ab[24][3] , \mult_23/ab[24][4] , \mult_23/ab[24][5] ,
         \mult_23/ab[24][6] , \mult_23/ab[24][7] , \mult_23/ab[25][0] ,
         \mult_23/ab[25][1] , \mult_23/ab[25][2] , \mult_23/ab[25][3] ,
         \mult_23/ab[25][4] , \mult_23/ab[25][5] , \mult_23/ab[25][6] ,
         \mult_23/ab[26][0] , \mult_23/ab[26][1] , \mult_23/ab[26][2] ,
         \mult_23/ab[26][3] , \mult_23/ab[26][4] , \mult_23/ab[26][5] ,
         \mult_23/ab[27][0] , \mult_23/ab[27][1] , \mult_23/ab[27][2] ,
         \mult_23/ab[27][3] , \mult_23/ab[27][4] , \mult_23/ab[28][0] ,
         \mult_23/ab[28][1] , \mult_23/ab[28][2] , \mult_23/ab[28][3] ,
         \mult_23/ab[29][0] , \mult_23/ab[29][1] , \mult_23/ab[29][2] ,
         \mult_23/ab[30][0] , \mult_23/ab[30][1] , \mult_23/ab[31][0] ;
  wire   [31:0] xy;
  wire   [31:0] o_reg;

  DFF \o_reg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[0])
         );
  DFF \o_reg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[1])
         );
  DFF \o_reg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[2])
         );
  DFF \o_reg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[3])
         );
  DFF \o_reg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[4])
         );
  DFF \o_reg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[5])
         );
  DFF \o_reg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[6])
         );
  DFF \o_reg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[7])
         );
  DFF \o_reg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[8])
         );
  DFF \o_reg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o_reg[9])
         );
  DFF \o_reg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[10]) );
  DFF \o_reg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[11]) );
  DFF \o_reg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[12]) );
  DFF \o_reg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[13]) );
  DFF \o_reg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[14]) );
  DFF \o_reg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[15]) );
  DFF \o_reg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[16]) );
  DFF \o_reg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[17]) );
  DFF \o_reg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[18]) );
  DFF \o_reg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[19]) );
  DFF \o_reg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[20]) );
  DFF \o_reg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[21]) );
  DFF \o_reg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[22]) );
  DFF \o_reg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[23]) );
  DFF \o_reg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[24]) );
  DFF \o_reg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[25]) );
  DFF \o_reg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[26]) );
  DFF \o_reg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[27]) );
  DFF \o_reg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[28]) );
  DFF \o_reg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[29]) );
  DFF \o_reg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[30]) );
  DFF \o_reg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        o_reg[31]) );
  FADDER \add_24/U1_1  ( .CIN(xy[1]), .IN0(o_reg[1]), .IN1(\add_24/carry[1] ), 
        .COUT(\add_24/carry[2] ), .SUM(o[1]) );
  FADDER \add_24/U1_2  ( .CIN(xy[2]), .IN0(o_reg[2]), .IN1(\add_24/carry[2] ), 
        .COUT(\add_24/carry[3] ), .SUM(o[2]) );
  FADDER \add_24/U1_3  ( .CIN(xy[3]), .IN0(o_reg[3]), .IN1(\add_24/carry[3] ), 
        .COUT(\add_24/carry[4] ), .SUM(o[3]) );
  FADDER \add_24/U1_4  ( .CIN(xy[4]), .IN0(o_reg[4]), .IN1(\add_24/carry[4] ), 
        .COUT(\add_24/carry[5] ), .SUM(o[4]) );
  FADDER \add_24/U1_5  ( .CIN(xy[5]), .IN0(o_reg[5]), .IN1(\add_24/carry[5] ), 
        .COUT(\add_24/carry[6] ), .SUM(o[5]) );
  FADDER \add_24/U1_6  ( .CIN(xy[6]), .IN0(o_reg[6]), .IN1(\add_24/carry[6] ), 
        .COUT(\add_24/carry[7] ), .SUM(o[6]) );
  FADDER \add_24/U1_7  ( .CIN(xy[7]), .IN0(o_reg[7]), .IN1(\add_24/carry[7] ), 
        .COUT(\add_24/carry[8] ), .SUM(o[7]) );
  FADDER \add_24/U1_8  ( .CIN(xy[8]), .IN0(o_reg[8]), .IN1(\add_24/carry[8] ), 
        .COUT(\add_24/carry[9] ), .SUM(o[8]) );
  FADDER \add_24/U1_9  ( .CIN(xy[9]), .IN0(o_reg[9]), .IN1(\add_24/carry[9] ), 
        .COUT(\add_24/carry[10] ), .SUM(o[9]) );
  FADDER \add_24/U1_10  ( .CIN(xy[10]), .IN0(o_reg[10]), .IN1(
        \add_24/carry[10] ), .COUT(\add_24/carry[11] ), .SUM(o[10]) );
  FADDER \add_24/U1_11  ( .CIN(xy[11]), .IN0(o_reg[11]), .IN1(
        \add_24/carry[11] ), .COUT(\add_24/carry[12] ), .SUM(o[11]) );
  FADDER \add_24/U1_12  ( .CIN(xy[12]), .IN0(o_reg[12]), .IN1(
        \add_24/carry[12] ), .COUT(\add_24/carry[13] ), .SUM(o[12]) );
  FADDER \add_24/U1_13  ( .CIN(xy[13]), .IN0(o_reg[13]), .IN1(
        \add_24/carry[13] ), .COUT(\add_24/carry[14] ), .SUM(o[13]) );
  FADDER \add_24/U1_14  ( .CIN(xy[14]), .IN0(o_reg[14]), .IN1(
        \add_24/carry[14] ), .COUT(\add_24/carry[15] ), .SUM(o[14]) );
  FADDER \add_24/U1_15  ( .CIN(xy[15]), .IN0(o_reg[15]), .IN1(
        \add_24/carry[15] ), .COUT(\add_24/carry[16] ), .SUM(o[15]) );
  FADDER \add_24/U1_16  ( .CIN(xy[16]), .IN0(o_reg[16]), .IN1(
        \add_24/carry[16] ), .COUT(\add_24/carry[17] ), .SUM(o[16]) );
  FADDER \add_24/U1_17  ( .CIN(xy[17]), .IN0(o_reg[17]), .IN1(
        \add_24/carry[17] ), .COUT(\add_24/carry[18] ), .SUM(o[17]) );
  FADDER \add_24/U1_18  ( .CIN(xy[18]), .IN0(o_reg[18]), .IN1(
        \add_24/carry[18] ), .COUT(\add_24/carry[19] ), .SUM(o[18]) );
  FADDER \add_24/U1_19  ( .CIN(xy[19]), .IN0(o_reg[19]), .IN1(
        \add_24/carry[19] ), .COUT(\add_24/carry[20] ), .SUM(o[19]) );
  FADDER \add_24/U1_20  ( .CIN(xy[20]), .IN0(o_reg[20]), .IN1(
        \add_24/carry[20] ), .COUT(\add_24/carry[21] ), .SUM(o[20]) );
  FADDER \add_24/U1_21  ( .CIN(xy[21]), .IN0(o_reg[21]), .IN1(
        \add_24/carry[21] ), .COUT(\add_24/carry[22] ), .SUM(o[21]) );
  FADDER \add_24/U1_22  ( .CIN(xy[22]), .IN0(o_reg[22]), .IN1(
        \add_24/carry[22] ), .COUT(\add_24/carry[23] ), .SUM(o[22]) );
  FADDER \add_24/U1_23  ( .CIN(xy[23]), .IN0(o_reg[23]), .IN1(
        \add_24/carry[23] ), .COUT(\add_24/carry[24] ), .SUM(o[23]) );
  FADDER \add_24/U1_24  ( .CIN(xy[24]), .IN0(o_reg[24]), .IN1(
        \add_24/carry[24] ), .COUT(\add_24/carry[25] ), .SUM(o[24]) );
  FADDER \add_24/U1_25  ( .CIN(xy[25]), .IN0(o_reg[25]), .IN1(
        \add_24/carry[25] ), .COUT(\add_24/carry[26] ), .SUM(o[25]) );
  FADDER \add_24/U1_26  ( .CIN(xy[26]), .IN0(o_reg[26]), .IN1(
        \add_24/carry[26] ), .COUT(\add_24/carry[27] ), .SUM(o[26]) );
  FADDER \add_24/U1_27  ( .CIN(xy[27]), .IN0(o_reg[27]), .IN1(
        \add_24/carry[27] ), .COUT(\add_24/carry[28] ), .SUM(o[27]) );
  FADDER \add_24/U1_28  ( .CIN(xy[28]), .IN0(o_reg[28]), .IN1(
        \add_24/carry[28] ), .COUT(\add_24/carry[29] ), .SUM(o[28]) );
  FADDER \add_24/U1_29  ( .CIN(xy[29]), .IN0(o_reg[29]), .IN1(
        \add_24/carry[29] ), .COUT(\add_24/carry[30] ), .SUM(o[29]) );
  FADDER \add_24/U1_30  ( .CIN(xy[30]), .IN0(o_reg[30]), .IN1(
        \add_24/carry[30] ), .COUT(\add_24/carry[31] ), .SUM(o[30]) );
  FADDER \add_24/U1_31  ( .CIN(\mult_23/SUMB[31][0] ), .IN0(o_reg[31]), .IN1(
        \add_24/carry[31] ), .SUM(o[31]) );
  FADDER \mult_23/S2_2_29  ( .CIN(\mult_23/ab[2][29] ), .IN0(
        \mult_23/CARRYB[1][29] ), .IN1(\mult_23/SUMB[1][30] ), .SUM(
        \mult_23/SUMB[2][29] ) );
  FADDER \mult_23/S2_2_28  ( .CIN(\mult_23/ab[2][28] ), .IN0(
        \mult_23/CARRYB[1][28] ), .IN1(\mult_23/SUMB[1][29] ), .COUT(
        \mult_23/CARRYB[2][28] ), .SUM(\mult_23/SUMB[2][28] ) );
  FADDER \mult_23/S2_2_27  ( .CIN(\mult_23/ab[2][27] ), .IN0(
        \mult_23/CARRYB[1][27] ), .IN1(\mult_23/SUMB[1][28] ), .COUT(
        \mult_23/CARRYB[2][27] ), .SUM(\mult_23/SUMB[2][27] ) );
  FADDER \mult_23/S2_2_26  ( .CIN(\mult_23/ab[2][26] ), .IN0(
        \mult_23/CARRYB[1][26] ), .IN1(\mult_23/SUMB[1][27] ), .COUT(
        \mult_23/CARRYB[2][26] ), .SUM(\mult_23/SUMB[2][26] ) );
  FADDER \mult_23/S2_2_25  ( .CIN(\mult_23/ab[2][25] ), .IN0(
        \mult_23/CARRYB[1][25] ), .IN1(\mult_23/SUMB[1][26] ), .COUT(
        \mult_23/CARRYB[2][25] ), .SUM(\mult_23/SUMB[2][25] ) );
  FADDER \mult_23/S2_2_24  ( .CIN(\mult_23/ab[2][24] ), .IN0(
        \mult_23/CARRYB[1][24] ), .IN1(\mult_23/SUMB[1][25] ), .COUT(
        \mult_23/CARRYB[2][24] ), .SUM(\mult_23/SUMB[2][24] ) );
  FADDER \mult_23/S2_2_23  ( .CIN(\mult_23/ab[2][23] ), .IN0(
        \mult_23/CARRYB[1][23] ), .IN1(\mult_23/SUMB[1][24] ), .COUT(
        \mult_23/CARRYB[2][23] ), .SUM(\mult_23/SUMB[2][23] ) );
  FADDER \mult_23/S2_2_22  ( .CIN(\mult_23/ab[2][22] ), .IN0(
        \mult_23/CARRYB[1][22] ), .IN1(\mult_23/SUMB[1][23] ), .COUT(
        \mult_23/CARRYB[2][22] ), .SUM(\mult_23/SUMB[2][22] ) );
  FADDER \mult_23/S2_2_21  ( .CIN(\mult_23/ab[2][21] ), .IN0(
        \mult_23/CARRYB[1][21] ), .IN1(\mult_23/SUMB[1][22] ), .COUT(
        \mult_23/CARRYB[2][21] ), .SUM(\mult_23/SUMB[2][21] ) );
  FADDER \mult_23/S2_2_20  ( .CIN(\mult_23/ab[2][20] ), .IN0(
        \mult_23/CARRYB[1][20] ), .IN1(\mult_23/SUMB[1][21] ), .COUT(
        \mult_23/CARRYB[2][20] ), .SUM(\mult_23/SUMB[2][20] ) );
  FADDER \mult_23/S2_2_19  ( .CIN(\mult_23/ab[2][19] ), .IN0(
        \mult_23/CARRYB[1][19] ), .IN1(\mult_23/SUMB[1][20] ), .COUT(
        \mult_23/CARRYB[2][19] ), .SUM(\mult_23/SUMB[2][19] ) );
  FADDER \mult_23/S2_2_18  ( .CIN(\mult_23/ab[2][18] ), .IN0(
        \mult_23/CARRYB[1][18] ), .IN1(\mult_23/SUMB[1][19] ), .COUT(
        \mult_23/CARRYB[2][18] ), .SUM(\mult_23/SUMB[2][18] ) );
  FADDER \mult_23/S2_2_17  ( .CIN(\mult_23/ab[2][17] ), .IN0(
        \mult_23/CARRYB[1][17] ), .IN1(\mult_23/SUMB[1][18] ), .COUT(
        \mult_23/CARRYB[2][17] ), .SUM(\mult_23/SUMB[2][17] ) );
  FADDER \mult_23/S2_2_16  ( .CIN(\mult_23/ab[2][16] ), .IN0(
        \mult_23/CARRYB[1][16] ), .IN1(\mult_23/SUMB[1][17] ), .COUT(
        \mult_23/CARRYB[2][16] ), .SUM(\mult_23/SUMB[2][16] ) );
  FADDER \mult_23/S2_2_15  ( .CIN(\mult_23/ab[2][15] ), .IN0(
        \mult_23/CARRYB[1][15] ), .IN1(\mult_23/SUMB[1][16] ), .COUT(
        \mult_23/CARRYB[2][15] ), .SUM(\mult_23/SUMB[2][15] ) );
  FADDER \mult_23/S2_2_14  ( .CIN(\mult_23/ab[2][14] ), .IN0(
        \mult_23/CARRYB[1][14] ), .IN1(\mult_23/SUMB[1][15] ), .COUT(
        \mult_23/CARRYB[2][14] ), .SUM(\mult_23/SUMB[2][14] ) );
  FADDER \mult_23/S2_2_13  ( .CIN(\mult_23/ab[2][13] ), .IN0(
        \mult_23/CARRYB[1][13] ), .IN1(\mult_23/SUMB[1][14] ), .COUT(
        \mult_23/CARRYB[2][13] ), .SUM(\mult_23/SUMB[2][13] ) );
  FADDER \mult_23/S2_2_12  ( .CIN(\mult_23/ab[2][12] ), .IN0(
        \mult_23/CARRYB[1][12] ), .IN1(\mult_23/SUMB[1][13] ), .COUT(
        \mult_23/CARRYB[2][12] ), .SUM(\mult_23/SUMB[2][12] ) );
  FADDER \mult_23/S2_2_11  ( .CIN(\mult_23/ab[2][11] ), .IN0(
        \mult_23/CARRYB[1][11] ), .IN1(\mult_23/SUMB[1][12] ), .COUT(
        \mult_23/CARRYB[2][11] ), .SUM(\mult_23/SUMB[2][11] ) );
  FADDER \mult_23/S2_2_10  ( .CIN(\mult_23/ab[2][10] ), .IN0(
        \mult_23/CARRYB[1][10] ), .IN1(\mult_23/SUMB[1][11] ), .COUT(
        \mult_23/CARRYB[2][10] ), .SUM(\mult_23/SUMB[2][10] ) );
  FADDER \mult_23/S2_2_9  ( .CIN(\mult_23/ab[2][9] ), .IN0(
        \mult_23/CARRYB[1][9] ), .IN1(\mult_23/SUMB[1][10] ), .COUT(
        \mult_23/CARRYB[2][9] ), .SUM(\mult_23/SUMB[2][9] ) );
  FADDER \mult_23/S2_2_8  ( .CIN(\mult_23/ab[2][8] ), .IN0(
        \mult_23/CARRYB[1][8] ), .IN1(\mult_23/SUMB[1][9] ), .COUT(
        \mult_23/CARRYB[2][8] ), .SUM(\mult_23/SUMB[2][8] ) );
  FADDER \mult_23/S2_2_7  ( .CIN(\mult_23/ab[2][7] ), .IN0(
        \mult_23/CARRYB[1][7] ), .IN1(\mult_23/SUMB[1][8] ), .COUT(
        \mult_23/CARRYB[2][7] ), .SUM(\mult_23/SUMB[2][7] ) );
  FADDER \mult_23/S2_2_6  ( .CIN(\mult_23/ab[2][6] ), .IN0(
        \mult_23/CARRYB[1][6] ), .IN1(\mult_23/SUMB[1][7] ), .COUT(
        \mult_23/CARRYB[2][6] ), .SUM(\mult_23/SUMB[2][6] ) );
  FADDER \mult_23/S2_2_5  ( .CIN(\mult_23/ab[2][5] ), .IN0(
        \mult_23/CARRYB[1][5] ), .IN1(\mult_23/SUMB[1][6] ), .COUT(
        \mult_23/CARRYB[2][5] ), .SUM(\mult_23/SUMB[2][5] ) );
  FADDER \mult_23/S2_2_4  ( .CIN(\mult_23/ab[2][4] ), .IN0(
        \mult_23/CARRYB[1][4] ), .IN1(\mult_23/SUMB[1][5] ), .COUT(
        \mult_23/CARRYB[2][4] ), .SUM(\mult_23/SUMB[2][4] ) );
  FADDER \mult_23/S2_2_3  ( .CIN(\mult_23/ab[2][3] ), .IN0(
        \mult_23/CARRYB[1][3] ), .IN1(\mult_23/SUMB[1][4] ), .COUT(
        \mult_23/CARRYB[2][3] ), .SUM(\mult_23/SUMB[2][3] ) );
  FADDER \mult_23/S2_2_2  ( .CIN(\mult_23/ab[2][2] ), .IN0(
        \mult_23/CARRYB[1][2] ), .IN1(\mult_23/SUMB[1][3] ), .COUT(
        \mult_23/CARRYB[2][2] ), .SUM(\mult_23/SUMB[2][2] ) );
  FADDER \mult_23/S2_2_1  ( .CIN(\mult_23/ab[2][1] ), .IN0(
        \mult_23/CARRYB[1][1] ), .IN1(\mult_23/SUMB[1][2] ), .COUT(
        \mult_23/CARRYB[2][1] ), .SUM(\mult_23/SUMB[2][1] ) );
  FADDER \mult_23/S1_2_0  ( .CIN(\mult_23/ab[2][0] ), .IN0(
        \mult_23/CARRYB[1][0] ), .IN1(\mult_23/SUMB[1][1] ), .COUT(
        \mult_23/CARRYB[2][0] ), .SUM(xy[2]) );
  FADDER \mult_23/S2_3_28  ( .CIN(\mult_23/ab[3][28] ), .IN0(
        \mult_23/CARRYB[2][28] ), .IN1(\mult_23/SUMB[2][29] ), .SUM(
        \mult_23/SUMB[3][28] ) );
  FADDER \mult_23/S2_3_27  ( .CIN(\mult_23/ab[3][27] ), .IN0(
        \mult_23/CARRYB[2][27] ), .IN1(\mult_23/SUMB[2][28] ), .COUT(
        \mult_23/CARRYB[3][27] ), .SUM(\mult_23/SUMB[3][27] ) );
  FADDER \mult_23/S2_3_26  ( .CIN(\mult_23/ab[3][26] ), .IN0(
        \mult_23/CARRYB[2][26] ), .IN1(\mult_23/SUMB[2][27] ), .COUT(
        \mult_23/CARRYB[3][26] ), .SUM(\mult_23/SUMB[3][26] ) );
  FADDER \mult_23/S2_3_25  ( .CIN(\mult_23/ab[3][25] ), .IN0(
        \mult_23/CARRYB[2][25] ), .IN1(\mult_23/SUMB[2][26] ), .COUT(
        \mult_23/CARRYB[3][25] ), .SUM(\mult_23/SUMB[3][25] ) );
  FADDER \mult_23/S2_3_24  ( .CIN(\mult_23/ab[3][24] ), .IN0(
        \mult_23/CARRYB[2][24] ), .IN1(\mult_23/SUMB[2][25] ), .COUT(
        \mult_23/CARRYB[3][24] ), .SUM(\mult_23/SUMB[3][24] ) );
  FADDER \mult_23/S2_3_23  ( .CIN(\mult_23/ab[3][23] ), .IN0(
        \mult_23/CARRYB[2][23] ), .IN1(\mult_23/SUMB[2][24] ), .COUT(
        \mult_23/CARRYB[3][23] ), .SUM(\mult_23/SUMB[3][23] ) );
  FADDER \mult_23/S2_3_22  ( .CIN(\mult_23/ab[3][22] ), .IN0(
        \mult_23/CARRYB[2][22] ), .IN1(\mult_23/SUMB[2][23] ), .COUT(
        \mult_23/CARRYB[3][22] ), .SUM(\mult_23/SUMB[3][22] ) );
  FADDER \mult_23/S2_3_21  ( .CIN(\mult_23/ab[3][21] ), .IN0(
        \mult_23/CARRYB[2][21] ), .IN1(\mult_23/SUMB[2][22] ), .COUT(
        \mult_23/CARRYB[3][21] ), .SUM(\mult_23/SUMB[3][21] ) );
  FADDER \mult_23/S2_3_20  ( .CIN(\mult_23/ab[3][20] ), .IN0(
        \mult_23/CARRYB[2][20] ), .IN1(\mult_23/SUMB[2][21] ), .COUT(
        \mult_23/CARRYB[3][20] ), .SUM(\mult_23/SUMB[3][20] ) );
  FADDER \mult_23/S2_3_19  ( .CIN(\mult_23/ab[3][19] ), .IN0(
        \mult_23/CARRYB[2][19] ), .IN1(\mult_23/SUMB[2][20] ), .COUT(
        \mult_23/CARRYB[3][19] ), .SUM(\mult_23/SUMB[3][19] ) );
  FADDER \mult_23/S2_3_18  ( .CIN(\mult_23/ab[3][18] ), .IN0(
        \mult_23/CARRYB[2][18] ), .IN1(\mult_23/SUMB[2][19] ), .COUT(
        \mult_23/CARRYB[3][18] ), .SUM(\mult_23/SUMB[3][18] ) );
  FADDER \mult_23/S2_3_17  ( .CIN(\mult_23/ab[3][17] ), .IN0(
        \mult_23/CARRYB[2][17] ), .IN1(\mult_23/SUMB[2][18] ), .COUT(
        \mult_23/CARRYB[3][17] ), .SUM(\mult_23/SUMB[3][17] ) );
  FADDER \mult_23/S2_3_16  ( .CIN(\mult_23/ab[3][16] ), .IN0(
        \mult_23/CARRYB[2][16] ), .IN1(\mult_23/SUMB[2][17] ), .COUT(
        \mult_23/CARRYB[3][16] ), .SUM(\mult_23/SUMB[3][16] ) );
  FADDER \mult_23/S2_3_15  ( .CIN(\mult_23/ab[3][15] ), .IN0(
        \mult_23/CARRYB[2][15] ), .IN1(\mult_23/SUMB[2][16] ), .COUT(
        \mult_23/CARRYB[3][15] ), .SUM(\mult_23/SUMB[3][15] ) );
  FADDER \mult_23/S2_3_14  ( .CIN(\mult_23/ab[3][14] ), .IN0(
        \mult_23/CARRYB[2][14] ), .IN1(\mult_23/SUMB[2][15] ), .COUT(
        \mult_23/CARRYB[3][14] ), .SUM(\mult_23/SUMB[3][14] ) );
  FADDER \mult_23/S2_3_13  ( .CIN(\mult_23/ab[3][13] ), .IN0(
        \mult_23/CARRYB[2][13] ), .IN1(\mult_23/SUMB[2][14] ), .COUT(
        \mult_23/CARRYB[3][13] ), .SUM(\mult_23/SUMB[3][13] ) );
  FADDER \mult_23/S2_3_12  ( .CIN(\mult_23/ab[3][12] ), .IN0(
        \mult_23/CARRYB[2][12] ), .IN1(\mult_23/SUMB[2][13] ), .COUT(
        \mult_23/CARRYB[3][12] ), .SUM(\mult_23/SUMB[3][12] ) );
  FADDER \mult_23/S2_3_11  ( .CIN(\mult_23/ab[3][11] ), .IN0(
        \mult_23/CARRYB[2][11] ), .IN1(\mult_23/SUMB[2][12] ), .COUT(
        \mult_23/CARRYB[3][11] ), .SUM(\mult_23/SUMB[3][11] ) );
  FADDER \mult_23/S2_3_10  ( .CIN(\mult_23/ab[3][10] ), .IN0(
        \mult_23/CARRYB[2][10] ), .IN1(\mult_23/SUMB[2][11] ), .COUT(
        \mult_23/CARRYB[3][10] ), .SUM(\mult_23/SUMB[3][10] ) );
  FADDER \mult_23/S2_3_9  ( .CIN(\mult_23/ab[3][9] ), .IN0(
        \mult_23/CARRYB[2][9] ), .IN1(\mult_23/SUMB[2][10] ), .COUT(
        \mult_23/CARRYB[3][9] ), .SUM(\mult_23/SUMB[3][9] ) );
  FADDER \mult_23/S2_3_8  ( .CIN(\mult_23/ab[3][8] ), .IN0(
        \mult_23/CARRYB[2][8] ), .IN1(\mult_23/SUMB[2][9] ), .COUT(
        \mult_23/CARRYB[3][8] ), .SUM(\mult_23/SUMB[3][8] ) );
  FADDER \mult_23/S2_3_7  ( .CIN(\mult_23/ab[3][7] ), .IN0(
        \mult_23/CARRYB[2][7] ), .IN1(\mult_23/SUMB[2][8] ), .COUT(
        \mult_23/CARRYB[3][7] ), .SUM(\mult_23/SUMB[3][7] ) );
  FADDER \mult_23/S2_3_6  ( .CIN(\mult_23/ab[3][6] ), .IN0(
        \mult_23/CARRYB[2][6] ), .IN1(\mult_23/SUMB[2][7] ), .COUT(
        \mult_23/CARRYB[3][6] ), .SUM(\mult_23/SUMB[3][6] ) );
  FADDER \mult_23/S2_3_5  ( .CIN(\mult_23/ab[3][5] ), .IN0(
        \mult_23/CARRYB[2][5] ), .IN1(\mult_23/SUMB[2][6] ), .COUT(
        \mult_23/CARRYB[3][5] ), .SUM(\mult_23/SUMB[3][5] ) );
  FADDER \mult_23/S2_3_4  ( .CIN(\mult_23/ab[3][4] ), .IN0(
        \mult_23/CARRYB[2][4] ), .IN1(\mult_23/SUMB[2][5] ), .COUT(
        \mult_23/CARRYB[3][4] ), .SUM(\mult_23/SUMB[3][4] ) );
  FADDER \mult_23/S2_3_3  ( .CIN(\mult_23/ab[3][3] ), .IN0(
        \mult_23/CARRYB[2][3] ), .IN1(\mult_23/SUMB[2][4] ), .COUT(
        \mult_23/CARRYB[3][3] ), .SUM(\mult_23/SUMB[3][3] ) );
  FADDER \mult_23/S2_3_2  ( .CIN(\mult_23/ab[3][2] ), .IN0(
        \mult_23/CARRYB[2][2] ), .IN1(\mult_23/SUMB[2][3] ), .COUT(
        \mult_23/CARRYB[3][2] ), .SUM(\mult_23/SUMB[3][2] ) );
  FADDER \mult_23/S2_3_1  ( .CIN(\mult_23/ab[3][1] ), .IN0(
        \mult_23/CARRYB[2][1] ), .IN1(\mult_23/SUMB[2][2] ), .COUT(
        \mult_23/CARRYB[3][1] ), .SUM(\mult_23/SUMB[3][1] ) );
  FADDER \mult_23/S1_3_0  ( .CIN(\mult_23/ab[3][0] ), .IN0(
        \mult_23/CARRYB[2][0] ), .IN1(\mult_23/SUMB[2][1] ), .COUT(
        \mult_23/CARRYB[3][0] ), .SUM(xy[3]) );
  FADDER \mult_23/S2_4_27  ( .CIN(\mult_23/ab[4][27] ), .IN0(
        \mult_23/CARRYB[3][27] ), .IN1(\mult_23/SUMB[3][28] ), .SUM(
        \mult_23/SUMB[4][27] ) );
  FADDER \mult_23/S2_4_26  ( .CIN(\mult_23/ab[4][26] ), .IN0(
        \mult_23/CARRYB[3][26] ), .IN1(\mult_23/SUMB[3][27] ), .COUT(
        \mult_23/CARRYB[4][26] ), .SUM(\mult_23/SUMB[4][26] ) );
  FADDER \mult_23/S2_4_25  ( .CIN(\mult_23/ab[4][25] ), .IN0(
        \mult_23/CARRYB[3][25] ), .IN1(\mult_23/SUMB[3][26] ), .COUT(
        \mult_23/CARRYB[4][25] ), .SUM(\mult_23/SUMB[4][25] ) );
  FADDER \mult_23/S2_4_24  ( .CIN(\mult_23/ab[4][24] ), .IN0(
        \mult_23/CARRYB[3][24] ), .IN1(\mult_23/SUMB[3][25] ), .COUT(
        \mult_23/CARRYB[4][24] ), .SUM(\mult_23/SUMB[4][24] ) );
  FADDER \mult_23/S2_4_23  ( .CIN(\mult_23/ab[4][23] ), .IN0(
        \mult_23/CARRYB[3][23] ), .IN1(\mult_23/SUMB[3][24] ), .COUT(
        \mult_23/CARRYB[4][23] ), .SUM(\mult_23/SUMB[4][23] ) );
  FADDER \mult_23/S2_4_22  ( .CIN(\mult_23/ab[4][22] ), .IN0(
        \mult_23/CARRYB[3][22] ), .IN1(\mult_23/SUMB[3][23] ), .COUT(
        \mult_23/CARRYB[4][22] ), .SUM(\mult_23/SUMB[4][22] ) );
  FADDER \mult_23/S2_4_21  ( .CIN(\mult_23/ab[4][21] ), .IN0(
        \mult_23/CARRYB[3][21] ), .IN1(\mult_23/SUMB[3][22] ), .COUT(
        \mult_23/CARRYB[4][21] ), .SUM(\mult_23/SUMB[4][21] ) );
  FADDER \mult_23/S2_4_20  ( .CIN(\mult_23/ab[4][20] ), .IN0(
        \mult_23/CARRYB[3][20] ), .IN1(\mult_23/SUMB[3][21] ), .COUT(
        \mult_23/CARRYB[4][20] ), .SUM(\mult_23/SUMB[4][20] ) );
  FADDER \mult_23/S2_4_19  ( .CIN(\mult_23/ab[4][19] ), .IN0(
        \mult_23/CARRYB[3][19] ), .IN1(\mult_23/SUMB[3][20] ), .COUT(
        \mult_23/CARRYB[4][19] ), .SUM(\mult_23/SUMB[4][19] ) );
  FADDER \mult_23/S2_4_18  ( .CIN(\mult_23/ab[4][18] ), .IN0(
        \mult_23/CARRYB[3][18] ), .IN1(\mult_23/SUMB[3][19] ), .COUT(
        \mult_23/CARRYB[4][18] ), .SUM(\mult_23/SUMB[4][18] ) );
  FADDER \mult_23/S2_4_17  ( .CIN(\mult_23/ab[4][17] ), .IN0(
        \mult_23/CARRYB[3][17] ), .IN1(\mult_23/SUMB[3][18] ), .COUT(
        \mult_23/CARRYB[4][17] ), .SUM(\mult_23/SUMB[4][17] ) );
  FADDER \mult_23/S2_4_16  ( .CIN(\mult_23/ab[4][16] ), .IN0(
        \mult_23/CARRYB[3][16] ), .IN1(\mult_23/SUMB[3][17] ), .COUT(
        \mult_23/CARRYB[4][16] ), .SUM(\mult_23/SUMB[4][16] ) );
  FADDER \mult_23/S2_4_15  ( .CIN(\mult_23/ab[4][15] ), .IN0(
        \mult_23/CARRYB[3][15] ), .IN1(\mult_23/SUMB[3][16] ), .COUT(
        \mult_23/CARRYB[4][15] ), .SUM(\mult_23/SUMB[4][15] ) );
  FADDER \mult_23/S2_4_14  ( .CIN(\mult_23/ab[4][14] ), .IN0(
        \mult_23/CARRYB[3][14] ), .IN1(\mult_23/SUMB[3][15] ), .COUT(
        \mult_23/CARRYB[4][14] ), .SUM(\mult_23/SUMB[4][14] ) );
  FADDER \mult_23/S2_4_13  ( .CIN(\mult_23/ab[4][13] ), .IN0(
        \mult_23/CARRYB[3][13] ), .IN1(\mult_23/SUMB[3][14] ), .COUT(
        \mult_23/CARRYB[4][13] ), .SUM(\mult_23/SUMB[4][13] ) );
  FADDER \mult_23/S2_4_12  ( .CIN(\mult_23/ab[4][12] ), .IN0(
        \mult_23/CARRYB[3][12] ), .IN1(\mult_23/SUMB[3][13] ), .COUT(
        \mult_23/CARRYB[4][12] ), .SUM(\mult_23/SUMB[4][12] ) );
  FADDER \mult_23/S2_4_11  ( .CIN(\mult_23/ab[4][11] ), .IN0(
        \mult_23/CARRYB[3][11] ), .IN1(\mult_23/SUMB[3][12] ), .COUT(
        \mult_23/CARRYB[4][11] ), .SUM(\mult_23/SUMB[4][11] ) );
  FADDER \mult_23/S2_4_10  ( .CIN(\mult_23/ab[4][10] ), .IN0(
        \mult_23/CARRYB[3][10] ), .IN1(\mult_23/SUMB[3][11] ), .COUT(
        \mult_23/CARRYB[4][10] ), .SUM(\mult_23/SUMB[4][10] ) );
  FADDER \mult_23/S2_4_9  ( .CIN(\mult_23/ab[4][9] ), .IN0(
        \mult_23/CARRYB[3][9] ), .IN1(\mult_23/SUMB[3][10] ), .COUT(
        \mult_23/CARRYB[4][9] ), .SUM(\mult_23/SUMB[4][9] ) );
  FADDER \mult_23/S2_4_8  ( .CIN(\mult_23/ab[4][8] ), .IN0(
        \mult_23/CARRYB[3][8] ), .IN1(\mult_23/SUMB[3][9] ), .COUT(
        \mult_23/CARRYB[4][8] ), .SUM(\mult_23/SUMB[4][8] ) );
  FADDER \mult_23/S2_4_7  ( .CIN(\mult_23/ab[4][7] ), .IN0(
        \mult_23/CARRYB[3][7] ), .IN1(\mult_23/SUMB[3][8] ), .COUT(
        \mult_23/CARRYB[4][7] ), .SUM(\mult_23/SUMB[4][7] ) );
  FADDER \mult_23/S2_4_6  ( .CIN(\mult_23/ab[4][6] ), .IN0(
        \mult_23/CARRYB[3][6] ), .IN1(\mult_23/SUMB[3][7] ), .COUT(
        \mult_23/CARRYB[4][6] ), .SUM(\mult_23/SUMB[4][6] ) );
  FADDER \mult_23/S2_4_5  ( .CIN(\mult_23/ab[4][5] ), .IN0(
        \mult_23/CARRYB[3][5] ), .IN1(\mult_23/SUMB[3][6] ), .COUT(
        \mult_23/CARRYB[4][5] ), .SUM(\mult_23/SUMB[4][5] ) );
  FADDER \mult_23/S2_4_4  ( .CIN(\mult_23/ab[4][4] ), .IN0(
        \mult_23/CARRYB[3][4] ), .IN1(\mult_23/SUMB[3][5] ), .COUT(
        \mult_23/CARRYB[4][4] ), .SUM(\mult_23/SUMB[4][4] ) );
  FADDER \mult_23/S2_4_3  ( .CIN(\mult_23/ab[4][3] ), .IN0(
        \mult_23/CARRYB[3][3] ), .IN1(\mult_23/SUMB[3][4] ), .COUT(
        \mult_23/CARRYB[4][3] ), .SUM(\mult_23/SUMB[4][3] ) );
  FADDER \mult_23/S2_4_2  ( .CIN(\mult_23/ab[4][2] ), .IN0(
        \mult_23/CARRYB[3][2] ), .IN1(\mult_23/SUMB[3][3] ), .COUT(
        \mult_23/CARRYB[4][2] ), .SUM(\mult_23/SUMB[4][2] ) );
  FADDER \mult_23/S2_4_1  ( .CIN(\mult_23/ab[4][1] ), .IN0(
        \mult_23/CARRYB[3][1] ), .IN1(\mult_23/SUMB[3][2] ), .COUT(
        \mult_23/CARRYB[4][1] ), .SUM(\mult_23/SUMB[4][1] ) );
  FADDER \mult_23/S1_4_0  ( .CIN(\mult_23/ab[4][0] ), .IN0(
        \mult_23/CARRYB[3][0] ), .IN1(\mult_23/SUMB[3][1] ), .COUT(
        \mult_23/CARRYB[4][0] ), .SUM(xy[4]) );
  FADDER \mult_23/S2_5_26  ( .CIN(\mult_23/ab[5][26] ), .IN0(
        \mult_23/CARRYB[4][26] ), .IN1(\mult_23/SUMB[4][27] ), .SUM(
        \mult_23/SUMB[5][26] ) );
  FADDER \mult_23/S2_5_25  ( .CIN(\mult_23/ab[5][25] ), .IN0(
        \mult_23/CARRYB[4][25] ), .IN1(\mult_23/SUMB[4][26] ), .COUT(
        \mult_23/CARRYB[5][25] ), .SUM(\mult_23/SUMB[5][25] ) );
  FADDER \mult_23/S2_5_24  ( .CIN(\mult_23/ab[5][24] ), .IN0(
        \mult_23/CARRYB[4][24] ), .IN1(\mult_23/SUMB[4][25] ), .COUT(
        \mult_23/CARRYB[5][24] ), .SUM(\mult_23/SUMB[5][24] ) );
  FADDER \mult_23/S2_5_23  ( .CIN(\mult_23/ab[5][23] ), .IN0(
        \mult_23/CARRYB[4][23] ), .IN1(\mult_23/SUMB[4][24] ), .COUT(
        \mult_23/CARRYB[5][23] ), .SUM(\mult_23/SUMB[5][23] ) );
  FADDER \mult_23/S2_5_22  ( .CIN(\mult_23/ab[5][22] ), .IN0(
        \mult_23/CARRYB[4][22] ), .IN1(\mult_23/SUMB[4][23] ), .COUT(
        \mult_23/CARRYB[5][22] ), .SUM(\mult_23/SUMB[5][22] ) );
  FADDER \mult_23/S2_5_21  ( .CIN(\mult_23/ab[5][21] ), .IN0(
        \mult_23/CARRYB[4][21] ), .IN1(\mult_23/SUMB[4][22] ), .COUT(
        \mult_23/CARRYB[5][21] ), .SUM(\mult_23/SUMB[5][21] ) );
  FADDER \mult_23/S2_5_20  ( .CIN(\mult_23/ab[5][20] ), .IN0(
        \mult_23/CARRYB[4][20] ), .IN1(\mult_23/SUMB[4][21] ), .COUT(
        \mult_23/CARRYB[5][20] ), .SUM(\mult_23/SUMB[5][20] ) );
  FADDER \mult_23/S2_5_19  ( .CIN(\mult_23/ab[5][19] ), .IN0(
        \mult_23/CARRYB[4][19] ), .IN1(\mult_23/SUMB[4][20] ), .COUT(
        \mult_23/CARRYB[5][19] ), .SUM(\mult_23/SUMB[5][19] ) );
  FADDER \mult_23/S2_5_18  ( .CIN(\mult_23/ab[5][18] ), .IN0(
        \mult_23/CARRYB[4][18] ), .IN1(\mult_23/SUMB[4][19] ), .COUT(
        \mult_23/CARRYB[5][18] ), .SUM(\mult_23/SUMB[5][18] ) );
  FADDER \mult_23/S2_5_17  ( .CIN(\mult_23/ab[5][17] ), .IN0(
        \mult_23/CARRYB[4][17] ), .IN1(\mult_23/SUMB[4][18] ), .COUT(
        \mult_23/CARRYB[5][17] ), .SUM(\mult_23/SUMB[5][17] ) );
  FADDER \mult_23/S2_5_16  ( .CIN(\mult_23/ab[5][16] ), .IN0(
        \mult_23/CARRYB[4][16] ), .IN1(\mult_23/SUMB[4][17] ), .COUT(
        \mult_23/CARRYB[5][16] ), .SUM(\mult_23/SUMB[5][16] ) );
  FADDER \mult_23/S2_5_15  ( .CIN(\mult_23/ab[5][15] ), .IN0(
        \mult_23/CARRYB[4][15] ), .IN1(\mult_23/SUMB[4][16] ), .COUT(
        \mult_23/CARRYB[5][15] ), .SUM(\mult_23/SUMB[5][15] ) );
  FADDER \mult_23/S2_5_14  ( .CIN(\mult_23/ab[5][14] ), .IN0(
        \mult_23/CARRYB[4][14] ), .IN1(\mult_23/SUMB[4][15] ), .COUT(
        \mult_23/CARRYB[5][14] ), .SUM(\mult_23/SUMB[5][14] ) );
  FADDER \mult_23/S2_5_13  ( .CIN(\mult_23/ab[5][13] ), .IN0(
        \mult_23/CARRYB[4][13] ), .IN1(\mult_23/SUMB[4][14] ), .COUT(
        \mult_23/CARRYB[5][13] ), .SUM(\mult_23/SUMB[5][13] ) );
  FADDER \mult_23/S2_5_12  ( .CIN(\mult_23/ab[5][12] ), .IN0(
        \mult_23/CARRYB[4][12] ), .IN1(\mult_23/SUMB[4][13] ), .COUT(
        \mult_23/CARRYB[5][12] ), .SUM(\mult_23/SUMB[5][12] ) );
  FADDER \mult_23/S2_5_11  ( .CIN(\mult_23/ab[5][11] ), .IN0(
        \mult_23/CARRYB[4][11] ), .IN1(\mult_23/SUMB[4][12] ), .COUT(
        \mult_23/CARRYB[5][11] ), .SUM(\mult_23/SUMB[5][11] ) );
  FADDER \mult_23/S2_5_10  ( .CIN(\mult_23/ab[5][10] ), .IN0(
        \mult_23/CARRYB[4][10] ), .IN1(\mult_23/SUMB[4][11] ), .COUT(
        \mult_23/CARRYB[5][10] ), .SUM(\mult_23/SUMB[5][10] ) );
  FADDER \mult_23/S2_5_9  ( .CIN(\mult_23/ab[5][9] ), .IN0(
        \mult_23/CARRYB[4][9] ), .IN1(\mult_23/SUMB[4][10] ), .COUT(
        \mult_23/CARRYB[5][9] ), .SUM(\mult_23/SUMB[5][9] ) );
  FADDER \mult_23/S2_5_8  ( .CIN(\mult_23/ab[5][8] ), .IN0(
        \mult_23/CARRYB[4][8] ), .IN1(\mult_23/SUMB[4][9] ), .COUT(
        \mult_23/CARRYB[5][8] ), .SUM(\mult_23/SUMB[5][8] ) );
  FADDER \mult_23/S2_5_7  ( .CIN(\mult_23/ab[5][7] ), .IN0(
        \mult_23/CARRYB[4][7] ), .IN1(\mult_23/SUMB[4][8] ), .COUT(
        \mult_23/CARRYB[5][7] ), .SUM(\mult_23/SUMB[5][7] ) );
  FADDER \mult_23/S2_5_6  ( .CIN(\mult_23/ab[5][6] ), .IN0(
        \mult_23/CARRYB[4][6] ), .IN1(\mult_23/SUMB[4][7] ), .COUT(
        \mult_23/CARRYB[5][6] ), .SUM(\mult_23/SUMB[5][6] ) );
  FADDER \mult_23/S2_5_5  ( .CIN(\mult_23/ab[5][5] ), .IN0(
        \mult_23/CARRYB[4][5] ), .IN1(\mult_23/SUMB[4][6] ), .COUT(
        \mult_23/CARRYB[5][5] ), .SUM(\mult_23/SUMB[5][5] ) );
  FADDER \mult_23/S2_5_4  ( .CIN(\mult_23/ab[5][4] ), .IN0(
        \mult_23/CARRYB[4][4] ), .IN1(\mult_23/SUMB[4][5] ), .COUT(
        \mult_23/CARRYB[5][4] ), .SUM(\mult_23/SUMB[5][4] ) );
  FADDER \mult_23/S2_5_3  ( .CIN(\mult_23/ab[5][3] ), .IN0(
        \mult_23/CARRYB[4][3] ), .IN1(\mult_23/SUMB[4][4] ), .COUT(
        \mult_23/CARRYB[5][3] ), .SUM(\mult_23/SUMB[5][3] ) );
  FADDER \mult_23/S2_5_2  ( .CIN(\mult_23/ab[5][2] ), .IN0(
        \mult_23/CARRYB[4][2] ), .IN1(\mult_23/SUMB[4][3] ), .COUT(
        \mult_23/CARRYB[5][2] ), .SUM(\mult_23/SUMB[5][2] ) );
  FADDER \mult_23/S2_5_1  ( .CIN(\mult_23/ab[5][1] ), .IN0(
        \mult_23/CARRYB[4][1] ), .IN1(\mult_23/SUMB[4][2] ), .COUT(
        \mult_23/CARRYB[5][1] ), .SUM(\mult_23/SUMB[5][1] ) );
  FADDER \mult_23/S1_5_0  ( .CIN(\mult_23/ab[5][0] ), .IN0(
        \mult_23/CARRYB[4][0] ), .IN1(\mult_23/SUMB[4][1] ), .COUT(
        \mult_23/CARRYB[5][0] ), .SUM(xy[5]) );
  FADDER \mult_23/S2_6_25  ( .CIN(\mult_23/ab[6][25] ), .IN0(
        \mult_23/CARRYB[5][25] ), .IN1(\mult_23/SUMB[5][26] ), .SUM(
        \mult_23/SUMB[6][25] ) );
  FADDER \mult_23/S2_6_24  ( .CIN(\mult_23/ab[6][24] ), .IN0(
        \mult_23/CARRYB[5][24] ), .IN1(\mult_23/SUMB[5][25] ), .COUT(
        \mult_23/CARRYB[6][24] ), .SUM(\mult_23/SUMB[6][24] ) );
  FADDER \mult_23/S2_6_23  ( .CIN(\mult_23/ab[6][23] ), .IN0(
        \mult_23/CARRYB[5][23] ), .IN1(\mult_23/SUMB[5][24] ), .COUT(
        \mult_23/CARRYB[6][23] ), .SUM(\mult_23/SUMB[6][23] ) );
  FADDER \mult_23/S2_6_22  ( .CIN(\mult_23/ab[6][22] ), .IN0(
        \mult_23/CARRYB[5][22] ), .IN1(\mult_23/SUMB[5][23] ), .COUT(
        \mult_23/CARRYB[6][22] ), .SUM(\mult_23/SUMB[6][22] ) );
  FADDER \mult_23/S2_6_21  ( .CIN(\mult_23/ab[6][21] ), .IN0(
        \mult_23/CARRYB[5][21] ), .IN1(\mult_23/SUMB[5][22] ), .COUT(
        \mult_23/CARRYB[6][21] ), .SUM(\mult_23/SUMB[6][21] ) );
  FADDER \mult_23/S2_6_20  ( .CIN(\mult_23/ab[6][20] ), .IN0(
        \mult_23/CARRYB[5][20] ), .IN1(\mult_23/SUMB[5][21] ), .COUT(
        \mult_23/CARRYB[6][20] ), .SUM(\mult_23/SUMB[6][20] ) );
  FADDER \mult_23/S2_6_19  ( .CIN(\mult_23/ab[6][19] ), .IN0(
        \mult_23/CARRYB[5][19] ), .IN1(\mult_23/SUMB[5][20] ), .COUT(
        \mult_23/CARRYB[6][19] ), .SUM(\mult_23/SUMB[6][19] ) );
  FADDER \mult_23/S2_6_18  ( .CIN(\mult_23/ab[6][18] ), .IN0(
        \mult_23/CARRYB[5][18] ), .IN1(\mult_23/SUMB[5][19] ), .COUT(
        \mult_23/CARRYB[6][18] ), .SUM(\mult_23/SUMB[6][18] ) );
  FADDER \mult_23/S2_6_17  ( .CIN(\mult_23/ab[6][17] ), .IN0(
        \mult_23/CARRYB[5][17] ), .IN1(\mult_23/SUMB[5][18] ), .COUT(
        \mult_23/CARRYB[6][17] ), .SUM(\mult_23/SUMB[6][17] ) );
  FADDER \mult_23/S2_6_16  ( .CIN(\mult_23/ab[6][16] ), .IN0(
        \mult_23/CARRYB[5][16] ), .IN1(\mult_23/SUMB[5][17] ), .COUT(
        \mult_23/CARRYB[6][16] ), .SUM(\mult_23/SUMB[6][16] ) );
  FADDER \mult_23/S2_6_15  ( .CIN(\mult_23/ab[6][15] ), .IN0(
        \mult_23/CARRYB[5][15] ), .IN1(\mult_23/SUMB[5][16] ), .COUT(
        \mult_23/CARRYB[6][15] ), .SUM(\mult_23/SUMB[6][15] ) );
  FADDER \mult_23/S2_6_14  ( .CIN(\mult_23/ab[6][14] ), .IN0(
        \mult_23/CARRYB[5][14] ), .IN1(\mult_23/SUMB[5][15] ), .COUT(
        \mult_23/CARRYB[6][14] ), .SUM(\mult_23/SUMB[6][14] ) );
  FADDER \mult_23/S2_6_13  ( .CIN(\mult_23/ab[6][13] ), .IN0(
        \mult_23/CARRYB[5][13] ), .IN1(\mult_23/SUMB[5][14] ), .COUT(
        \mult_23/CARRYB[6][13] ), .SUM(\mult_23/SUMB[6][13] ) );
  FADDER \mult_23/S2_6_12  ( .CIN(\mult_23/ab[6][12] ), .IN0(
        \mult_23/CARRYB[5][12] ), .IN1(\mult_23/SUMB[5][13] ), .COUT(
        \mult_23/CARRYB[6][12] ), .SUM(\mult_23/SUMB[6][12] ) );
  FADDER \mult_23/S2_6_11  ( .CIN(\mult_23/ab[6][11] ), .IN0(
        \mult_23/CARRYB[5][11] ), .IN1(\mult_23/SUMB[5][12] ), .COUT(
        \mult_23/CARRYB[6][11] ), .SUM(\mult_23/SUMB[6][11] ) );
  FADDER \mult_23/S2_6_10  ( .CIN(\mult_23/ab[6][10] ), .IN0(
        \mult_23/CARRYB[5][10] ), .IN1(\mult_23/SUMB[5][11] ), .COUT(
        \mult_23/CARRYB[6][10] ), .SUM(\mult_23/SUMB[6][10] ) );
  FADDER \mult_23/S2_6_9  ( .CIN(\mult_23/ab[6][9] ), .IN0(
        \mult_23/CARRYB[5][9] ), .IN1(\mult_23/SUMB[5][10] ), .COUT(
        \mult_23/CARRYB[6][9] ), .SUM(\mult_23/SUMB[6][9] ) );
  FADDER \mult_23/S2_6_8  ( .CIN(\mult_23/ab[6][8] ), .IN0(
        \mult_23/CARRYB[5][8] ), .IN1(\mult_23/SUMB[5][9] ), .COUT(
        \mult_23/CARRYB[6][8] ), .SUM(\mult_23/SUMB[6][8] ) );
  FADDER \mult_23/S2_6_7  ( .CIN(\mult_23/ab[6][7] ), .IN0(
        \mult_23/CARRYB[5][7] ), .IN1(\mult_23/SUMB[5][8] ), .COUT(
        \mult_23/CARRYB[6][7] ), .SUM(\mult_23/SUMB[6][7] ) );
  FADDER \mult_23/S2_6_6  ( .CIN(\mult_23/ab[6][6] ), .IN0(
        \mult_23/CARRYB[5][6] ), .IN1(\mult_23/SUMB[5][7] ), .COUT(
        \mult_23/CARRYB[6][6] ), .SUM(\mult_23/SUMB[6][6] ) );
  FADDER \mult_23/S2_6_5  ( .CIN(\mult_23/ab[6][5] ), .IN0(
        \mult_23/CARRYB[5][5] ), .IN1(\mult_23/SUMB[5][6] ), .COUT(
        \mult_23/CARRYB[6][5] ), .SUM(\mult_23/SUMB[6][5] ) );
  FADDER \mult_23/S2_6_4  ( .CIN(\mult_23/ab[6][4] ), .IN0(
        \mult_23/CARRYB[5][4] ), .IN1(\mult_23/SUMB[5][5] ), .COUT(
        \mult_23/CARRYB[6][4] ), .SUM(\mult_23/SUMB[6][4] ) );
  FADDER \mult_23/S2_6_3  ( .CIN(\mult_23/ab[6][3] ), .IN0(
        \mult_23/CARRYB[5][3] ), .IN1(\mult_23/SUMB[5][4] ), .COUT(
        \mult_23/CARRYB[6][3] ), .SUM(\mult_23/SUMB[6][3] ) );
  FADDER \mult_23/S2_6_2  ( .CIN(\mult_23/ab[6][2] ), .IN0(
        \mult_23/CARRYB[5][2] ), .IN1(\mult_23/SUMB[5][3] ), .COUT(
        \mult_23/CARRYB[6][2] ), .SUM(\mult_23/SUMB[6][2] ) );
  FADDER \mult_23/S2_6_1  ( .CIN(\mult_23/ab[6][1] ), .IN0(
        \mult_23/CARRYB[5][1] ), .IN1(\mult_23/SUMB[5][2] ), .COUT(
        \mult_23/CARRYB[6][1] ), .SUM(\mult_23/SUMB[6][1] ) );
  FADDER \mult_23/S1_6_0  ( .CIN(\mult_23/ab[6][0] ), .IN0(
        \mult_23/CARRYB[5][0] ), .IN1(\mult_23/SUMB[5][1] ), .COUT(
        \mult_23/CARRYB[6][0] ), .SUM(xy[6]) );
  FADDER \mult_23/S2_7_24  ( .CIN(\mult_23/ab[7][24] ), .IN0(
        \mult_23/CARRYB[6][24] ), .IN1(\mult_23/SUMB[6][25] ), .SUM(
        \mult_23/SUMB[7][24] ) );
  FADDER \mult_23/S2_7_23  ( .CIN(\mult_23/ab[7][23] ), .IN0(
        \mult_23/CARRYB[6][23] ), .IN1(\mult_23/SUMB[6][24] ), .COUT(
        \mult_23/CARRYB[7][23] ), .SUM(\mult_23/SUMB[7][23] ) );
  FADDER \mult_23/S2_7_22  ( .CIN(\mult_23/ab[7][22] ), .IN0(
        \mult_23/CARRYB[6][22] ), .IN1(\mult_23/SUMB[6][23] ), .COUT(
        \mult_23/CARRYB[7][22] ), .SUM(\mult_23/SUMB[7][22] ) );
  FADDER \mult_23/S2_7_21  ( .CIN(\mult_23/ab[7][21] ), .IN0(
        \mult_23/CARRYB[6][21] ), .IN1(\mult_23/SUMB[6][22] ), .COUT(
        \mult_23/CARRYB[7][21] ), .SUM(\mult_23/SUMB[7][21] ) );
  FADDER \mult_23/S2_7_20  ( .CIN(\mult_23/ab[7][20] ), .IN0(
        \mult_23/CARRYB[6][20] ), .IN1(\mult_23/SUMB[6][21] ), .COUT(
        \mult_23/CARRYB[7][20] ), .SUM(\mult_23/SUMB[7][20] ) );
  FADDER \mult_23/S2_7_19  ( .CIN(\mult_23/ab[7][19] ), .IN0(
        \mult_23/CARRYB[6][19] ), .IN1(\mult_23/SUMB[6][20] ), .COUT(
        \mult_23/CARRYB[7][19] ), .SUM(\mult_23/SUMB[7][19] ) );
  FADDER \mult_23/S2_7_18  ( .CIN(\mult_23/ab[7][18] ), .IN0(
        \mult_23/CARRYB[6][18] ), .IN1(\mult_23/SUMB[6][19] ), .COUT(
        \mult_23/CARRYB[7][18] ), .SUM(\mult_23/SUMB[7][18] ) );
  FADDER \mult_23/S2_7_17  ( .CIN(\mult_23/ab[7][17] ), .IN0(
        \mult_23/CARRYB[6][17] ), .IN1(\mult_23/SUMB[6][18] ), .COUT(
        \mult_23/CARRYB[7][17] ), .SUM(\mult_23/SUMB[7][17] ) );
  FADDER \mult_23/S2_7_16  ( .CIN(\mult_23/ab[7][16] ), .IN0(
        \mult_23/CARRYB[6][16] ), .IN1(\mult_23/SUMB[6][17] ), .COUT(
        \mult_23/CARRYB[7][16] ), .SUM(\mult_23/SUMB[7][16] ) );
  FADDER \mult_23/S2_7_15  ( .CIN(\mult_23/ab[7][15] ), .IN0(
        \mult_23/CARRYB[6][15] ), .IN1(\mult_23/SUMB[6][16] ), .COUT(
        \mult_23/CARRYB[7][15] ), .SUM(\mult_23/SUMB[7][15] ) );
  FADDER \mult_23/S2_7_14  ( .CIN(\mult_23/ab[7][14] ), .IN0(
        \mult_23/CARRYB[6][14] ), .IN1(\mult_23/SUMB[6][15] ), .COUT(
        \mult_23/CARRYB[7][14] ), .SUM(\mult_23/SUMB[7][14] ) );
  FADDER \mult_23/S2_7_13  ( .CIN(\mult_23/ab[7][13] ), .IN0(
        \mult_23/CARRYB[6][13] ), .IN1(\mult_23/SUMB[6][14] ), .COUT(
        \mult_23/CARRYB[7][13] ), .SUM(\mult_23/SUMB[7][13] ) );
  FADDER \mult_23/S2_7_12  ( .CIN(\mult_23/ab[7][12] ), .IN0(
        \mult_23/CARRYB[6][12] ), .IN1(\mult_23/SUMB[6][13] ), .COUT(
        \mult_23/CARRYB[7][12] ), .SUM(\mult_23/SUMB[7][12] ) );
  FADDER \mult_23/S2_7_11  ( .CIN(\mult_23/ab[7][11] ), .IN0(
        \mult_23/CARRYB[6][11] ), .IN1(\mult_23/SUMB[6][12] ), .COUT(
        \mult_23/CARRYB[7][11] ), .SUM(\mult_23/SUMB[7][11] ) );
  FADDER \mult_23/S2_7_10  ( .CIN(\mult_23/ab[7][10] ), .IN0(
        \mult_23/CARRYB[6][10] ), .IN1(\mult_23/SUMB[6][11] ), .COUT(
        \mult_23/CARRYB[7][10] ), .SUM(\mult_23/SUMB[7][10] ) );
  FADDER \mult_23/S2_7_9  ( .CIN(\mult_23/ab[7][9] ), .IN0(
        \mult_23/CARRYB[6][9] ), .IN1(\mult_23/SUMB[6][10] ), .COUT(
        \mult_23/CARRYB[7][9] ), .SUM(\mult_23/SUMB[7][9] ) );
  FADDER \mult_23/S2_7_8  ( .CIN(\mult_23/ab[7][8] ), .IN0(
        \mult_23/CARRYB[6][8] ), .IN1(\mult_23/SUMB[6][9] ), .COUT(
        \mult_23/CARRYB[7][8] ), .SUM(\mult_23/SUMB[7][8] ) );
  FADDER \mult_23/S2_7_7  ( .CIN(\mult_23/ab[7][7] ), .IN0(
        \mult_23/CARRYB[6][7] ), .IN1(\mult_23/SUMB[6][8] ), .COUT(
        \mult_23/CARRYB[7][7] ), .SUM(\mult_23/SUMB[7][7] ) );
  FADDER \mult_23/S2_7_6  ( .CIN(\mult_23/ab[7][6] ), .IN0(
        \mult_23/CARRYB[6][6] ), .IN1(\mult_23/SUMB[6][7] ), .COUT(
        \mult_23/CARRYB[7][6] ), .SUM(\mult_23/SUMB[7][6] ) );
  FADDER \mult_23/S2_7_5  ( .CIN(\mult_23/ab[7][5] ), .IN0(
        \mult_23/CARRYB[6][5] ), .IN1(\mult_23/SUMB[6][6] ), .COUT(
        \mult_23/CARRYB[7][5] ), .SUM(\mult_23/SUMB[7][5] ) );
  FADDER \mult_23/S2_7_4  ( .CIN(\mult_23/ab[7][4] ), .IN0(
        \mult_23/CARRYB[6][4] ), .IN1(\mult_23/SUMB[6][5] ), .COUT(
        \mult_23/CARRYB[7][4] ), .SUM(\mult_23/SUMB[7][4] ) );
  FADDER \mult_23/S2_7_3  ( .CIN(\mult_23/ab[7][3] ), .IN0(
        \mult_23/CARRYB[6][3] ), .IN1(\mult_23/SUMB[6][4] ), .COUT(
        \mult_23/CARRYB[7][3] ), .SUM(\mult_23/SUMB[7][3] ) );
  FADDER \mult_23/S2_7_2  ( .CIN(\mult_23/ab[7][2] ), .IN0(
        \mult_23/CARRYB[6][2] ), .IN1(\mult_23/SUMB[6][3] ), .COUT(
        \mult_23/CARRYB[7][2] ), .SUM(\mult_23/SUMB[7][2] ) );
  FADDER \mult_23/S2_7_1  ( .CIN(\mult_23/ab[7][1] ), .IN0(
        \mult_23/CARRYB[6][1] ), .IN1(\mult_23/SUMB[6][2] ), .COUT(
        \mult_23/CARRYB[7][1] ), .SUM(\mult_23/SUMB[7][1] ) );
  FADDER \mult_23/S1_7_0  ( .CIN(\mult_23/ab[7][0] ), .IN0(
        \mult_23/CARRYB[6][0] ), .IN1(\mult_23/SUMB[6][1] ), .COUT(
        \mult_23/CARRYB[7][0] ), .SUM(xy[7]) );
  FADDER \mult_23/S2_8_23  ( .CIN(\mult_23/ab[8][23] ), .IN0(
        \mult_23/CARRYB[7][23] ), .IN1(\mult_23/SUMB[7][24] ), .SUM(
        \mult_23/SUMB[8][23] ) );
  FADDER \mult_23/S2_8_22  ( .CIN(\mult_23/ab[8][22] ), .IN0(
        \mult_23/CARRYB[7][22] ), .IN1(\mult_23/SUMB[7][23] ), .COUT(
        \mult_23/CARRYB[8][22] ), .SUM(\mult_23/SUMB[8][22] ) );
  FADDER \mult_23/S2_8_21  ( .CIN(\mult_23/ab[8][21] ), .IN0(
        \mult_23/CARRYB[7][21] ), .IN1(\mult_23/SUMB[7][22] ), .COUT(
        \mult_23/CARRYB[8][21] ), .SUM(\mult_23/SUMB[8][21] ) );
  FADDER \mult_23/S2_8_20  ( .CIN(\mult_23/ab[8][20] ), .IN0(
        \mult_23/CARRYB[7][20] ), .IN1(\mult_23/SUMB[7][21] ), .COUT(
        \mult_23/CARRYB[8][20] ), .SUM(\mult_23/SUMB[8][20] ) );
  FADDER \mult_23/S2_8_19  ( .CIN(\mult_23/ab[8][19] ), .IN0(
        \mult_23/CARRYB[7][19] ), .IN1(\mult_23/SUMB[7][20] ), .COUT(
        \mult_23/CARRYB[8][19] ), .SUM(\mult_23/SUMB[8][19] ) );
  FADDER \mult_23/S2_8_18  ( .CIN(\mult_23/ab[8][18] ), .IN0(
        \mult_23/CARRYB[7][18] ), .IN1(\mult_23/SUMB[7][19] ), .COUT(
        \mult_23/CARRYB[8][18] ), .SUM(\mult_23/SUMB[8][18] ) );
  FADDER \mult_23/S2_8_17  ( .CIN(\mult_23/ab[8][17] ), .IN0(
        \mult_23/CARRYB[7][17] ), .IN1(\mult_23/SUMB[7][18] ), .COUT(
        \mult_23/CARRYB[8][17] ), .SUM(\mult_23/SUMB[8][17] ) );
  FADDER \mult_23/S2_8_16  ( .CIN(\mult_23/ab[8][16] ), .IN0(
        \mult_23/CARRYB[7][16] ), .IN1(\mult_23/SUMB[7][17] ), .COUT(
        \mult_23/CARRYB[8][16] ), .SUM(\mult_23/SUMB[8][16] ) );
  FADDER \mult_23/S2_8_15  ( .CIN(\mult_23/ab[8][15] ), .IN0(
        \mult_23/CARRYB[7][15] ), .IN1(\mult_23/SUMB[7][16] ), .COUT(
        \mult_23/CARRYB[8][15] ), .SUM(\mult_23/SUMB[8][15] ) );
  FADDER \mult_23/S2_8_14  ( .CIN(\mult_23/ab[8][14] ), .IN0(
        \mult_23/CARRYB[7][14] ), .IN1(\mult_23/SUMB[7][15] ), .COUT(
        \mult_23/CARRYB[8][14] ), .SUM(\mult_23/SUMB[8][14] ) );
  FADDER \mult_23/S2_8_13  ( .CIN(\mult_23/ab[8][13] ), .IN0(
        \mult_23/CARRYB[7][13] ), .IN1(\mult_23/SUMB[7][14] ), .COUT(
        \mult_23/CARRYB[8][13] ), .SUM(\mult_23/SUMB[8][13] ) );
  FADDER \mult_23/S2_8_12  ( .CIN(\mult_23/ab[8][12] ), .IN0(
        \mult_23/CARRYB[7][12] ), .IN1(\mult_23/SUMB[7][13] ), .COUT(
        \mult_23/CARRYB[8][12] ), .SUM(\mult_23/SUMB[8][12] ) );
  FADDER \mult_23/S2_8_11  ( .CIN(\mult_23/ab[8][11] ), .IN0(
        \mult_23/CARRYB[7][11] ), .IN1(\mult_23/SUMB[7][12] ), .COUT(
        \mult_23/CARRYB[8][11] ), .SUM(\mult_23/SUMB[8][11] ) );
  FADDER \mult_23/S2_8_10  ( .CIN(\mult_23/ab[8][10] ), .IN0(
        \mult_23/CARRYB[7][10] ), .IN1(\mult_23/SUMB[7][11] ), .COUT(
        \mult_23/CARRYB[8][10] ), .SUM(\mult_23/SUMB[8][10] ) );
  FADDER \mult_23/S2_8_9  ( .CIN(\mult_23/ab[8][9] ), .IN0(
        \mult_23/CARRYB[7][9] ), .IN1(\mult_23/SUMB[7][10] ), .COUT(
        \mult_23/CARRYB[8][9] ), .SUM(\mult_23/SUMB[8][9] ) );
  FADDER \mult_23/S2_8_8  ( .CIN(\mult_23/ab[8][8] ), .IN0(
        \mult_23/CARRYB[7][8] ), .IN1(\mult_23/SUMB[7][9] ), .COUT(
        \mult_23/CARRYB[8][8] ), .SUM(\mult_23/SUMB[8][8] ) );
  FADDER \mult_23/S2_8_7  ( .CIN(\mult_23/ab[8][7] ), .IN0(
        \mult_23/CARRYB[7][7] ), .IN1(\mult_23/SUMB[7][8] ), .COUT(
        \mult_23/CARRYB[8][7] ), .SUM(\mult_23/SUMB[8][7] ) );
  FADDER \mult_23/S2_8_6  ( .CIN(\mult_23/ab[8][6] ), .IN0(
        \mult_23/CARRYB[7][6] ), .IN1(\mult_23/SUMB[7][7] ), .COUT(
        \mult_23/CARRYB[8][6] ), .SUM(\mult_23/SUMB[8][6] ) );
  FADDER \mult_23/S2_8_5  ( .CIN(\mult_23/ab[8][5] ), .IN0(
        \mult_23/CARRYB[7][5] ), .IN1(\mult_23/SUMB[7][6] ), .COUT(
        \mult_23/CARRYB[8][5] ), .SUM(\mult_23/SUMB[8][5] ) );
  FADDER \mult_23/S2_8_4  ( .CIN(\mult_23/ab[8][4] ), .IN0(
        \mult_23/CARRYB[7][4] ), .IN1(\mult_23/SUMB[7][5] ), .COUT(
        \mult_23/CARRYB[8][4] ), .SUM(\mult_23/SUMB[8][4] ) );
  FADDER \mult_23/S2_8_3  ( .CIN(\mult_23/ab[8][3] ), .IN0(
        \mult_23/CARRYB[7][3] ), .IN1(\mult_23/SUMB[7][4] ), .COUT(
        \mult_23/CARRYB[8][3] ), .SUM(\mult_23/SUMB[8][3] ) );
  FADDER \mult_23/S2_8_2  ( .CIN(\mult_23/ab[8][2] ), .IN0(
        \mult_23/CARRYB[7][2] ), .IN1(\mult_23/SUMB[7][3] ), .COUT(
        \mult_23/CARRYB[8][2] ), .SUM(\mult_23/SUMB[8][2] ) );
  FADDER \mult_23/S2_8_1  ( .CIN(\mult_23/ab[8][1] ), .IN0(
        \mult_23/CARRYB[7][1] ), .IN1(\mult_23/SUMB[7][2] ), .COUT(
        \mult_23/CARRYB[8][1] ), .SUM(\mult_23/SUMB[8][1] ) );
  FADDER \mult_23/S1_8_0  ( .CIN(\mult_23/ab[8][0] ), .IN0(
        \mult_23/CARRYB[7][0] ), .IN1(\mult_23/SUMB[7][1] ), .COUT(
        \mult_23/CARRYB[8][0] ), .SUM(xy[8]) );
  FADDER \mult_23/S2_9_22  ( .CIN(\mult_23/ab[9][22] ), .IN0(
        \mult_23/CARRYB[8][22] ), .IN1(\mult_23/SUMB[8][23] ), .SUM(
        \mult_23/SUMB[9][22] ) );
  FADDER \mult_23/S2_9_21  ( .CIN(\mult_23/ab[9][21] ), .IN0(
        \mult_23/CARRYB[8][21] ), .IN1(\mult_23/SUMB[8][22] ), .COUT(
        \mult_23/CARRYB[9][21] ), .SUM(\mult_23/SUMB[9][21] ) );
  FADDER \mult_23/S2_9_20  ( .CIN(\mult_23/ab[9][20] ), .IN0(
        \mult_23/CARRYB[8][20] ), .IN1(\mult_23/SUMB[8][21] ), .COUT(
        \mult_23/CARRYB[9][20] ), .SUM(\mult_23/SUMB[9][20] ) );
  FADDER \mult_23/S2_9_19  ( .CIN(\mult_23/ab[9][19] ), .IN0(
        \mult_23/CARRYB[8][19] ), .IN1(\mult_23/SUMB[8][20] ), .COUT(
        \mult_23/CARRYB[9][19] ), .SUM(\mult_23/SUMB[9][19] ) );
  FADDER \mult_23/S2_9_18  ( .CIN(\mult_23/ab[9][18] ), .IN0(
        \mult_23/CARRYB[8][18] ), .IN1(\mult_23/SUMB[8][19] ), .COUT(
        \mult_23/CARRYB[9][18] ), .SUM(\mult_23/SUMB[9][18] ) );
  FADDER \mult_23/S2_9_17  ( .CIN(\mult_23/ab[9][17] ), .IN0(
        \mult_23/CARRYB[8][17] ), .IN1(\mult_23/SUMB[8][18] ), .COUT(
        \mult_23/CARRYB[9][17] ), .SUM(\mult_23/SUMB[9][17] ) );
  FADDER \mult_23/S2_9_16  ( .CIN(\mult_23/ab[9][16] ), .IN0(
        \mult_23/CARRYB[8][16] ), .IN1(\mult_23/SUMB[8][17] ), .COUT(
        \mult_23/CARRYB[9][16] ), .SUM(\mult_23/SUMB[9][16] ) );
  FADDER \mult_23/S2_9_15  ( .CIN(\mult_23/ab[9][15] ), .IN0(
        \mult_23/CARRYB[8][15] ), .IN1(\mult_23/SUMB[8][16] ), .COUT(
        \mult_23/CARRYB[9][15] ), .SUM(\mult_23/SUMB[9][15] ) );
  FADDER \mult_23/S2_9_14  ( .CIN(\mult_23/ab[9][14] ), .IN0(
        \mult_23/CARRYB[8][14] ), .IN1(\mult_23/SUMB[8][15] ), .COUT(
        \mult_23/CARRYB[9][14] ), .SUM(\mult_23/SUMB[9][14] ) );
  FADDER \mult_23/S2_9_13  ( .CIN(\mult_23/ab[9][13] ), .IN0(
        \mult_23/CARRYB[8][13] ), .IN1(\mult_23/SUMB[8][14] ), .COUT(
        \mult_23/CARRYB[9][13] ), .SUM(\mult_23/SUMB[9][13] ) );
  FADDER \mult_23/S2_9_12  ( .CIN(\mult_23/ab[9][12] ), .IN0(
        \mult_23/CARRYB[8][12] ), .IN1(\mult_23/SUMB[8][13] ), .COUT(
        \mult_23/CARRYB[9][12] ), .SUM(\mult_23/SUMB[9][12] ) );
  FADDER \mult_23/S2_9_11  ( .CIN(\mult_23/ab[9][11] ), .IN0(
        \mult_23/CARRYB[8][11] ), .IN1(\mult_23/SUMB[8][12] ), .COUT(
        \mult_23/CARRYB[9][11] ), .SUM(\mult_23/SUMB[9][11] ) );
  FADDER \mult_23/S2_9_10  ( .CIN(\mult_23/ab[9][10] ), .IN0(
        \mult_23/CARRYB[8][10] ), .IN1(\mult_23/SUMB[8][11] ), .COUT(
        \mult_23/CARRYB[9][10] ), .SUM(\mult_23/SUMB[9][10] ) );
  FADDER \mult_23/S2_9_9  ( .CIN(\mult_23/ab[9][9] ), .IN0(
        \mult_23/CARRYB[8][9] ), .IN1(\mult_23/SUMB[8][10] ), .COUT(
        \mult_23/CARRYB[9][9] ), .SUM(\mult_23/SUMB[9][9] ) );
  FADDER \mult_23/S2_9_8  ( .CIN(\mult_23/ab[9][8] ), .IN0(
        \mult_23/CARRYB[8][8] ), .IN1(\mult_23/SUMB[8][9] ), .COUT(
        \mult_23/CARRYB[9][8] ), .SUM(\mult_23/SUMB[9][8] ) );
  FADDER \mult_23/S2_9_7  ( .CIN(\mult_23/ab[9][7] ), .IN0(
        \mult_23/CARRYB[8][7] ), .IN1(\mult_23/SUMB[8][8] ), .COUT(
        \mult_23/CARRYB[9][7] ), .SUM(\mult_23/SUMB[9][7] ) );
  FADDER \mult_23/S2_9_6  ( .CIN(\mult_23/ab[9][6] ), .IN0(
        \mult_23/CARRYB[8][6] ), .IN1(\mult_23/SUMB[8][7] ), .COUT(
        \mult_23/CARRYB[9][6] ), .SUM(\mult_23/SUMB[9][6] ) );
  FADDER \mult_23/S2_9_5  ( .CIN(\mult_23/ab[9][5] ), .IN0(
        \mult_23/CARRYB[8][5] ), .IN1(\mult_23/SUMB[8][6] ), .COUT(
        \mult_23/CARRYB[9][5] ), .SUM(\mult_23/SUMB[9][5] ) );
  FADDER \mult_23/S2_9_4  ( .CIN(\mult_23/ab[9][4] ), .IN0(
        \mult_23/CARRYB[8][4] ), .IN1(\mult_23/SUMB[8][5] ), .COUT(
        \mult_23/CARRYB[9][4] ), .SUM(\mult_23/SUMB[9][4] ) );
  FADDER \mult_23/S2_9_3  ( .CIN(\mult_23/ab[9][3] ), .IN0(
        \mult_23/CARRYB[8][3] ), .IN1(\mult_23/SUMB[8][4] ), .COUT(
        \mult_23/CARRYB[9][3] ), .SUM(\mult_23/SUMB[9][3] ) );
  FADDER \mult_23/S2_9_2  ( .CIN(\mult_23/ab[9][2] ), .IN0(
        \mult_23/CARRYB[8][2] ), .IN1(\mult_23/SUMB[8][3] ), .COUT(
        \mult_23/CARRYB[9][2] ), .SUM(\mult_23/SUMB[9][2] ) );
  FADDER \mult_23/S2_9_1  ( .CIN(\mult_23/ab[9][1] ), .IN0(
        \mult_23/CARRYB[8][1] ), .IN1(\mult_23/SUMB[8][2] ), .COUT(
        \mult_23/CARRYB[9][1] ), .SUM(\mult_23/SUMB[9][1] ) );
  FADDER \mult_23/S1_9_0  ( .CIN(\mult_23/ab[9][0] ), .IN0(
        \mult_23/CARRYB[8][0] ), .IN1(\mult_23/SUMB[8][1] ), .COUT(
        \mult_23/CARRYB[9][0] ), .SUM(xy[9]) );
  FADDER \mult_23/S2_10_21  ( .CIN(\mult_23/ab[10][21] ), .IN0(
        \mult_23/CARRYB[9][21] ), .IN1(\mult_23/SUMB[9][22] ), .SUM(
        \mult_23/SUMB[10][21] ) );
  FADDER \mult_23/S2_10_20  ( .CIN(\mult_23/ab[10][20] ), .IN0(
        \mult_23/CARRYB[9][20] ), .IN1(\mult_23/SUMB[9][21] ), .COUT(
        \mult_23/CARRYB[10][20] ), .SUM(\mult_23/SUMB[10][20] ) );
  FADDER \mult_23/S2_10_19  ( .CIN(\mult_23/ab[10][19] ), .IN0(
        \mult_23/CARRYB[9][19] ), .IN1(\mult_23/SUMB[9][20] ), .COUT(
        \mult_23/CARRYB[10][19] ), .SUM(\mult_23/SUMB[10][19] ) );
  FADDER \mult_23/S2_10_18  ( .CIN(\mult_23/ab[10][18] ), .IN0(
        \mult_23/CARRYB[9][18] ), .IN1(\mult_23/SUMB[9][19] ), .COUT(
        \mult_23/CARRYB[10][18] ), .SUM(\mult_23/SUMB[10][18] ) );
  FADDER \mult_23/S2_10_17  ( .CIN(\mult_23/ab[10][17] ), .IN0(
        \mult_23/CARRYB[9][17] ), .IN1(\mult_23/SUMB[9][18] ), .COUT(
        \mult_23/CARRYB[10][17] ), .SUM(\mult_23/SUMB[10][17] ) );
  FADDER \mult_23/S2_10_16  ( .CIN(\mult_23/ab[10][16] ), .IN0(
        \mult_23/CARRYB[9][16] ), .IN1(\mult_23/SUMB[9][17] ), .COUT(
        \mult_23/CARRYB[10][16] ), .SUM(\mult_23/SUMB[10][16] ) );
  FADDER \mult_23/S2_10_15  ( .CIN(\mult_23/ab[10][15] ), .IN0(
        \mult_23/CARRYB[9][15] ), .IN1(\mult_23/SUMB[9][16] ), .COUT(
        \mult_23/CARRYB[10][15] ), .SUM(\mult_23/SUMB[10][15] ) );
  FADDER \mult_23/S2_10_14  ( .CIN(\mult_23/ab[10][14] ), .IN0(
        \mult_23/CARRYB[9][14] ), .IN1(\mult_23/SUMB[9][15] ), .COUT(
        \mult_23/CARRYB[10][14] ), .SUM(\mult_23/SUMB[10][14] ) );
  FADDER \mult_23/S2_10_13  ( .CIN(\mult_23/ab[10][13] ), .IN0(
        \mult_23/CARRYB[9][13] ), .IN1(\mult_23/SUMB[9][14] ), .COUT(
        \mult_23/CARRYB[10][13] ), .SUM(\mult_23/SUMB[10][13] ) );
  FADDER \mult_23/S2_10_12  ( .CIN(\mult_23/ab[10][12] ), .IN0(
        \mult_23/CARRYB[9][12] ), .IN1(\mult_23/SUMB[9][13] ), .COUT(
        \mult_23/CARRYB[10][12] ), .SUM(\mult_23/SUMB[10][12] ) );
  FADDER \mult_23/S2_10_11  ( .CIN(\mult_23/ab[10][11] ), .IN0(
        \mult_23/CARRYB[9][11] ), .IN1(\mult_23/SUMB[9][12] ), .COUT(
        \mult_23/CARRYB[10][11] ), .SUM(\mult_23/SUMB[10][11] ) );
  FADDER \mult_23/S2_10_10  ( .CIN(\mult_23/ab[10][10] ), .IN0(
        \mult_23/CARRYB[9][10] ), .IN1(\mult_23/SUMB[9][11] ), .COUT(
        \mult_23/CARRYB[10][10] ), .SUM(\mult_23/SUMB[10][10] ) );
  FADDER \mult_23/S2_10_9  ( .CIN(\mult_23/ab[10][9] ), .IN0(
        \mult_23/CARRYB[9][9] ), .IN1(\mult_23/SUMB[9][10] ), .COUT(
        \mult_23/CARRYB[10][9] ), .SUM(\mult_23/SUMB[10][9] ) );
  FADDER \mult_23/S2_10_8  ( .CIN(\mult_23/ab[10][8] ), .IN0(
        \mult_23/CARRYB[9][8] ), .IN1(\mult_23/SUMB[9][9] ), .COUT(
        \mult_23/CARRYB[10][8] ), .SUM(\mult_23/SUMB[10][8] ) );
  FADDER \mult_23/S2_10_7  ( .CIN(\mult_23/ab[10][7] ), .IN0(
        \mult_23/CARRYB[9][7] ), .IN1(\mult_23/SUMB[9][8] ), .COUT(
        \mult_23/CARRYB[10][7] ), .SUM(\mult_23/SUMB[10][7] ) );
  FADDER \mult_23/S2_10_6  ( .CIN(\mult_23/ab[10][6] ), .IN0(
        \mult_23/CARRYB[9][6] ), .IN1(\mult_23/SUMB[9][7] ), .COUT(
        \mult_23/CARRYB[10][6] ), .SUM(\mult_23/SUMB[10][6] ) );
  FADDER \mult_23/S2_10_5  ( .CIN(\mult_23/ab[10][5] ), .IN0(
        \mult_23/CARRYB[9][5] ), .IN1(\mult_23/SUMB[9][6] ), .COUT(
        \mult_23/CARRYB[10][5] ), .SUM(\mult_23/SUMB[10][5] ) );
  FADDER \mult_23/S2_10_4  ( .CIN(\mult_23/ab[10][4] ), .IN0(
        \mult_23/CARRYB[9][4] ), .IN1(\mult_23/SUMB[9][5] ), .COUT(
        \mult_23/CARRYB[10][4] ), .SUM(\mult_23/SUMB[10][4] ) );
  FADDER \mult_23/S2_10_3  ( .CIN(\mult_23/ab[10][3] ), .IN0(
        \mult_23/CARRYB[9][3] ), .IN1(\mult_23/SUMB[9][4] ), .COUT(
        \mult_23/CARRYB[10][3] ), .SUM(\mult_23/SUMB[10][3] ) );
  FADDER \mult_23/S2_10_2  ( .CIN(\mult_23/ab[10][2] ), .IN0(
        \mult_23/CARRYB[9][2] ), .IN1(\mult_23/SUMB[9][3] ), .COUT(
        \mult_23/CARRYB[10][2] ), .SUM(\mult_23/SUMB[10][2] ) );
  FADDER \mult_23/S2_10_1  ( .CIN(\mult_23/ab[10][1] ), .IN0(
        \mult_23/CARRYB[9][1] ), .IN1(\mult_23/SUMB[9][2] ), .COUT(
        \mult_23/CARRYB[10][1] ), .SUM(\mult_23/SUMB[10][1] ) );
  FADDER \mult_23/S1_10_0  ( .CIN(\mult_23/ab[10][0] ), .IN0(
        \mult_23/CARRYB[9][0] ), .IN1(\mult_23/SUMB[9][1] ), .COUT(
        \mult_23/CARRYB[10][0] ), .SUM(xy[10]) );
  FADDER \mult_23/S2_11_20  ( .CIN(\mult_23/ab[11][20] ), .IN0(
        \mult_23/CARRYB[10][20] ), .IN1(\mult_23/SUMB[10][21] ), .SUM(
        \mult_23/SUMB[11][20] ) );
  FADDER \mult_23/S2_11_19  ( .CIN(\mult_23/ab[11][19] ), .IN0(
        \mult_23/CARRYB[10][19] ), .IN1(\mult_23/SUMB[10][20] ), .COUT(
        \mult_23/CARRYB[11][19] ), .SUM(\mult_23/SUMB[11][19] ) );
  FADDER \mult_23/S2_11_18  ( .CIN(\mult_23/ab[11][18] ), .IN0(
        \mult_23/CARRYB[10][18] ), .IN1(\mult_23/SUMB[10][19] ), .COUT(
        \mult_23/CARRYB[11][18] ), .SUM(\mult_23/SUMB[11][18] ) );
  FADDER \mult_23/S2_11_17  ( .CIN(\mult_23/ab[11][17] ), .IN0(
        \mult_23/CARRYB[10][17] ), .IN1(\mult_23/SUMB[10][18] ), .COUT(
        \mult_23/CARRYB[11][17] ), .SUM(\mult_23/SUMB[11][17] ) );
  FADDER \mult_23/S2_11_16  ( .CIN(\mult_23/ab[11][16] ), .IN0(
        \mult_23/CARRYB[10][16] ), .IN1(\mult_23/SUMB[10][17] ), .COUT(
        \mult_23/CARRYB[11][16] ), .SUM(\mult_23/SUMB[11][16] ) );
  FADDER \mult_23/S2_11_15  ( .CIN(\mult_23/ab[11][15] ), .IN0(
        \mult_23/CARRYB[10][15] ), .IN1(\mult_23/SUMB[10][16] ), .COUT(
        \mult_23/CARRYB[11][15] ), .SUM(\mult_23/SUMB[11][15] ) );
  FADDER \mult_23/S2_11_14  ( .CIN(\mult_23/ab[11][14] ), .IN0(
        \mult_23/CARRYB[10][14] ), .IN1(\mult_23/SUMB[10][15] ), .COUT(
        \mult_23/CARRYB[11][14] ), .SUM(\mult_23/SUMB[11][14] ) );
  FADDER \mult_23/S2_11_13  ( .CIN(\mult_23/ab[11][13] ), .IN0(
        \mult_23/CARRYB[10][13] ), .IN1(\mult_23/SUMB[10][14] ), .COUT(
        \mult_23/CARRYB[11][13] ), .SUM(\mult_23/SUMB[11][13] ) );
  FADDER \mult_23/S2_11_12  ( .CIN(\mult_23/ab[11][12] ), .IN0(
        \mult_23/CARRYB[10][12] ), .IN1(\mult_23/SUMB[10][13] ), .COUT(
        \mult_23/CARRYB[11][12] ), .SUM(\mult_23/SUMB[11][12] ) );
  FADDER \mult_23/S2_11_11  ( .CIN(\mult_23/ab[11][11] ), .IN0(
        \mult_23/CARRYB[10][11] ), .IN1(\mult_23/SUMB[10][12] ), .COUT(
        \mult_23/CARRYB[11][11] ), .SUM(\mult_23/SUMB[11][11] ) );
  FADDER \mult_23/S2_11_10  ( .CIN(\mult_23/ab[11][10] ), .IN0(
        \mult_23/CARRYB[10][10] ), .IN1(\mult_23/SUMB[10][11] ), .COUT(
        \mult_23/CARRYB[11][10] ), .SUM(\mult_23/SUMB[11][10] ) );
  FADDER \mult_23/S2_11_9  ( .CIN(\mult_23/ab[11][9] ), .IN0(
        \mult_23/CARRYB[10][9] ), .IN1(\mult_23/SUMB[10][10] ), .COUT(
        \mult_23/CARRYB[11][9] ), .SUM(\mult_23/SUMB[11][9] ) );
  FADDER \mult_23/S2_11_8  ( .CIN(\mult_23/ab[11][8] ), .IN0(
        \mult_23/CARRYB[10][8] ), .IN1(\mult_23/SUMB[10][9] ), .COUT(
        \mult_23/CARRYB[11][8] ), .SUM(\mult_23/SUMB[11][8] ) );
  FADDER \mult_23/S2_11_7  ( .CIN(\mult_23/ab[11][7] ), .IN0(
        \mult_23/CARRYB[10][7] ), .IN1(\mult_23/SUMB[10][8] ), .COUT(
        \mult_23/CARRYB[11][7] ), .SUM(\mult_23/SUMB[11][7] ) );
  FADDER \mult_23/S2_11_6  ( .CIN(\mult_23/ab[11][6] ), .IN0(
        \mult_23/CARRYB[10][6] ), .IN1(\mult_23/SUMB[10][7] ), .COUT(
        \mult_23/CARRYB[11][6] ), .SUM(\mult_23/SUMB[11][6] ) );
  FADDER \mult_23/S2_11_5  ( .CIN(\mult_23/ab[11][5] ), .IN0(
        \mult_23/CARRYB[10][5] ), .IN1(\mult_23/SUMB[10][6] ), .COUT(
        \mult_23/CARRYB[11][5] ), .SUM(\mult_23/SUMB[11][5] ) );
  FADDER \mult_23/S2_11_4  ( .CIN(\mult_23/ab[11][4] ), .IN0(
        \mult_23/CARRYB[10][4] ), .IN1(\mult_23/SUMB[10][5] ), .COUT(
        \mult_23/CARRYB[11][4] ), .SUM(\mult_23/SUMB[11][4] ) );
  FADDER \mult_23/S2_11_3  ( .CIN(\mult_23/ab[11][3] ), .IN0(
        \mult_23/CARRYB[10][3] ), .IN1(\mult_23/SUMB[10][4] ), .COUT(
        \mult_23/CARRYB[11][3] ), .SUM(\mult_23/SUMB[11][3] ) );
  FADDER \mult_23/S2_11_2  ( .CIN(\mult_23/ab[11][2] ), .IN0(
        \mult_23/CARRYB[10][2] ), .IN1(\mult_23/SUMB[10][3] ), .COUT(
        \mult_23/CARRYB[11][2] ), .SUM(\mult_23/SUMB[11][2] ) );
  FADDER \mult_23/S2_11_1  ( .CIN(\mult_23/ab[11][1] ), .IN0(
        \mult_23/CARRYB[10][1] ), .IN1(\mult_23/SUMB[10][2] ), .COUT(
        \mult_23/CARRYB[11][1] ), .SUM(\mult_23/SUMB[11][1] ) );
  FADDER \mult_23/S1_11_0  ( .CIN(\mult_23/ab[11][0] ), .IN0(
        \mult_23/CARRYB[10][0] ), .IN1(\mult_23/SUMB[10][1] ), .COUT(
        \mult_23/CARRYB[11][0] ), .SUM(xy[11]) );
  FADDER \mult_23/S2_12_19  ( .CIN(\mult_23/ab[12][19] ), .IN0(
        \mult_23/CARRYB[11][19] ), .IN1(\mult_23/SUMB[11][20] ), .SUM(
        \mult_23/SUMB[12][19] ) );
  FADDER \mult_23/S2_12_18  ( .CIN(\mult_23/ab[12][18] ), .IN0(
        \mult_23/CARRYB[11][18] ), .IN1(\mult_23/SUMB[11][19] ), .COUT(
        \mult_23/CARRYB[12][18] ), .SUM(\mult_23/SUMB[12][18] ) );
  FADDER \mult_23/S2_12_17  ( .CIN(\mult_23/ab[12][17] ), .IN0(
        \mult_23/CARRYB[11][17] ), .IN1(\mult_23/SUMB[11][18] ), .COUT(
        \mult_23/CARRYB[12][17] ), .SUM(\mult_23/SUMB[12][17] ) );
  FADDER \mult_23/S2_12_16  ( .CIN(\mult_23/ab[12][16] ), .IN0(
        \mult_23/CARRYB[11][16] ), .IN1(\mult_23/SUMB[11][17] ), .COUT(
        \mult_23/CARRYB[12][16] ), .SUM(\mult_23/SUMB[12][16] ) );
  FADDER \mult_23/S2_12_15  ( .CIN(\mult_23/ab[12][15] ), .IN0(
        \mult_23/CARRYB[11][15] ), .IN1(\mult_23/SUMB[11][16] ), .COUT(
        \mult_23/CARRYB[12][15] ), .SUM(\mult_23/SUMB[12][15] ) );
  FADDER \mult_23/S2_12_14  ( .CIN(\mult_23/ab[12][14] ), .IN0(
        \mult_23/CARRYB[11][14] ), .IN1(\mult_23/SUMB[11][15] ), .COUT(
        \mult_23/CARRYB[12][14] ), .SUM(\mult_23/SUMB[12][14] ) );
  FADDER \mult_23/S2_12_13  ( .CIN(\mult_23/ab[12][13] ), .IN0(
        \mult_23/CARRYB[11][13] ), .IN1(\mult_23/SUMB[11][14] ), .COUT(
        \mult_23/CARRYB[12][13] ), .SUM(\mult_23/SUMB[12][13] ) );
  FADDER \mult_23/S2_12_12  ( .CIN(\mult_23/ab[12][12] ), .IN0(
        \mult_23/CARRYB[11][12] ), .IN1(\mult_23/SUMB[11][13] ), .COUT(
        \mult_23/CARRYB[12][12] ), .SUM(\mult_23/SUMB[12][12] ) );
  FADDER \mult_23/S2_12_11  ( .CIN(\mult_23/ab[12][11] ), .IN0(
        \mult_23/CARRYB[11][11] ), .IN1(\mult_23/SUMB[11][12] ), .COUT(
        \mult_23/CARRYB[12][11] ), .SUM(\mult_23/SUMB[12][11] ) );
  FADDER \mult_23/S2_12_10  ( .CIN(\mult_23/ab[12][10] ), .IN0(
        \mult_23/CARRYB[11][10] ), .IN1(\mult_23/SUMB[11][11] ), .COUT(
        \mult_23/CARRYB[12][10] ), .SUM(\mult_23/SUMB[12][10] ) );
  FADDER \mult_23/S2_12_9  ( .CIN(\mult_23/ab[12][9] ), .IN0(
        \mult_23/CARRYB[11][9] ), .IN1(\mult_23/SUMB[11][10] ), .COUT(
        \mult_23/CARRYB[12][9] ), .SUM(\mult_23/SUMB[12][9] ) );
  FADDER \mult_23/S2_12_8  ( .CIN(\mult_23/ab[12][8] ), .IN0(
        \mult_23/CARRYB[11][8] ), .IN1(\mult_23/SUMB[11][9] ), .COUT(
        \mult_23/CARRYB[12][8] ), .SUM(\mult_23/SUMB[12][8] ) );
  FADDER \mult_23/S2_12_7  ( .CIN(\mult_23/ab[12][7] ), .IN0(
        \mult_23/CARRYB[11][7] ), .IN1(\mult_23/SUMB[11][8] ), .COUT(
        \mult_23/CARRYB[12][7] ), .SUM(\mult_23/SUMB[12][7] ) );
  FADDER \mult_23/S2_12_6  ( .CIN(\mult_23/ab[12][6] ), .IN0(
        \mult_23/CARRYB[11][6] ), .IN1(\mult_23/SUMB[11][7] ), .COUT(
        \mult_23/CARRYB[12][6] ), .SUM(\mult_23/SUMB[12][6] ) );
  FADDER \mult_23/S2_12_5  ( .CIN(\mult_23/ab[12][5] ), .IN0(
        \mult_23/CARRYB[11][5] ), .IN1(\mult_23/SUMB[11][6] ), .COUT(
        \mult_23/CARRYB[12][5] ), .SUM(\mult_23/SUMB[12][5] ) );
  FADDER \mult_23/S2_12_4  ( .CIN(\mult_23/ab[12][4] ), .IN0(
        \mult_23/CARRYB[11][4] ), .IN1(\mult_23/SUMB[11][5] ), .COUT(
        \mult_23/CARRYB[12][4] ), .SUM(\mult_23/SUMB[12][4] ) );
  FADDER \mult_23/S2_12_3  ( .CIN(\mult_23/ab[12][3] ), .IN0(
        \mult_23/CARRYB[11][3] ), .IN1(\mult_23/SUMB[11][4] ), .COUT(
        \mult_23/CARRYB[12][3] ), .SUM(\mult_23/SUMB[12][3] ) );
  FADDER \mult_23/S2_12_2  ( .CIN(\mult_23/ab[12][2] ), .IN0(
        \mult_23/CARRYB[11][2] ), .IN1(\mult_23/SUMB[11][3] ), .COUT(
        \mult_23/CARRYB[12][2] ), .SUM(\mult_23/SUMB[12][2] ) );
  FADDER \mult_23/S2_12_1  ( .CIN(\mult_23/ab[12][1] ), .IN0(
        \mult_23/CARRYB[11][1] ), .IN1(\mult_23/SUMB[11][2] ), .COUT(
        \mult_23/CARRYB[12][1] ), .SUM(\mult_23/SUMB[12][1] ) );
  FADDER \mult_23/S1_12_0  ( .CIN(\mult_23/ab[12][0] ), .IN0(
        \mult_23/CARRYB[11][0] ), .IN1(\mult_23/SUMB[11][1] ), .COUT(
        \mult_23/CARRYB[12][0] ), .SUM(xy[12]) );
  FADDER \mult_23/S2_13_18  ( .CIN(\mult_23/ab[13][18] ), .IN0(
        \mult_23/CARRYB[12][18] ), .IN1(\mult_23/SUMB[12][19] ), .SUM(
        \mult_23/SUMB[13][18] ) );
  FADDER \mult_23/S2_13_17  ( .CIN(\mult_23/ab[13][17] ), .IN0(
        \mult_23/CARRYB[12][17] ), .IN1(\mult_23/SUMB[12][18] ), .COUT(
        \mult_23/CARRYB[13][17] ), .SUM(\mult_23/SUMB[13][17] ) );
  FADDER \mult_23/S2_13_16  ( .CIN(\mult_23/ab[13][16] ), .IN0(
        \mult_23/CARRYB[12][16] ), .IN1(\mult_23/SUMB[12][17] ), .COUT(
        \mult_23/CARRYB[13][16] ), .SUM(\mult_23/SUMB[13][16] ) );
  FADDER \mult_23/S2_13_15  ( .CIN(\mult_23/ab[13][15] ), .IN0(
        \mult_23/CARRYB[12][15] ), .IN1(\mult_23/SUMB[12][16] ), .COUT(
        \mult_23/CARRYB[13][15] ), .SUM(\mult_23/SUMB[13][15] ) );
  FADDER \mult_23/S2_13_14  ( .CIN(\mult_23/ab[13][14] ), .IN0(
        \mult_23/CARRYB[12][14] ), .IN1(\mult_23/SUMB[12][15] ), .COUT(
        \mult_23/CARRYB[13][14] ), .SUM(\mult_23/SUMB[13][14] ) );
  FADDER \mult_23/S2_13_13  ( .CIN(\mult_23/ab[13][13] ), .IN0(
        \mult_23/CARRYB[12][13] ), .IN1(\mult_23/SUMB[12][14] ), .COUT(
        \mult_23/CARRYB[13][13] ), .SUM(\mult_23/SUMB[13][13] ) );
  FADDER \mult_23/S2_13_12  ( .CIN(\mult_23/ab[13][12] ), .IN0(
        \mult_23/CARRYB[12][12] ), .IN1(\mult_23/SUMB[12][13] ), .COUT(
        \mult_23/CARRYB[13][12] ), .SUM(\mult_23/SUMB[13][12] ) );
  FADDER \mult_23/S2_13_11  ( .CIN(\mult_23/ab[13][11] ), .IN0(
        \mult_23/CARRYB[12][11] ), .IN1(\mult_23/SUMB[12][12] ), .COUT(
        \mult_23/CARRYB[13][11] ), .SUM(\mult_23/SUMB[13][11] ) );
  FADDER \mult_23/S2_13_10  ( .CIN(\mult_23/ab[13][10] ), .IN0(
        \mult_23/CARRYB[12][10] ), .IN1(\mult_23/SUMB[12][11] ), .COUT(
        \mult_23/CARRYB[13][10] ), .SUM(\mult_23/SUMB[13][10] ) );
  FADDER \mult_23/S2_13_9  ( .CIN(\mult_23/ab[13][9] ), .IN0(
        \mult_23/CARRYB[12][9] ), .IN1(\mult_23/SUMB[12][10] ), .COUT(
        \mult_23/CARRYB[13][9] ), .SUM(\mult_23/SUMB[13][9] ) );
  FADDER \mult_23/S2_13_8  ( .CIN(\mult_23/ab[13][8] ), .IN0(
        \mult_23/CARRYB[12][8] ), .IN1(\mult_23/SUMB[12][9] ), .COUT(
        \mult_23/CARRYB[13][8] ), .SUM(\mult_23/SUMB[13][8] ) );
  FADDER \mult_23/S2_13_7  ( .CIN(\mult_23/ab[13][7] ), .IN0(
        \mult_23/CARRYB[12][7] ), .IN1(\mult_23/SUMB[12][8] ), .COUT(
        \mult_23/CARRYB[13][7] ), .SUM(\mult_23/SUMB[13][7] ) );
  FADDER \mult_23/S2_13_6  ( .CIN(\mult_23/ab[13][6] ), .IN0(
        \mult_23/CARRYB[12][6] ), .IN1(\mult_23/SUMB[12][7] ), .COUT(
        \mult_23/CARRYB[13][6] ), .SUM(\mult_23/SUMB[13][6] ) );
  FADDER \mult_23/S2_13_5  ( .CIN(\mult_23/ab[13][5] ), .IN0(
        \mult_23/CARRYB[12][5] ), .IN1(\mult_23/SUMB[12][6] ), .COUT(
        \mult_23/CARRYB[13][5] ), .SUM(\mult_23/SUMB[13][5] ) );
  FADDER \mult_23/S2_13_4  ( .CIN(\mult_23/ab[13][4] ), .IN0(
        \mult_23/CARRYB[12][4] ), .IN1(\mult_23/SUMB[12][5] ), .COUT(
        \mult_23/CARRYB[13][4] ), .SUM(\mult_23/SUMB[13][4] ) );
  FADDER \mult_23/S2_13_3  ( .CIN(\mult_23/ab[13][3] ), .IN0(
        \mult_23/CARRYB[12][3] ), .IN1(\mult_23/SUMB[12][4] ), .COUT(
        \mult_23/CARRYB[13][3] ), .SUM(\mult_23/SUMB[13][3] ) );
  FADDER \mult_23/S2_13_2  ( .CIN(\mult_23/ab[13][2] ), .IN0(
        \mult_23/CARRYB[12][2] ), .IN1(\mult_23/SUMB[12][3] ), .COUT(
        \mult_23/CARRYB[13][2] ), .SUM(\mult_23/SUMB[13][2] ) );
  FADDER \mult_23/S2_13_1  ( .CIN(\mult_23/ab[13][1] ), .IN0(
        \mult_23/CARRYB[12][1] ), .IN1(\mult_23/SUMB[12][2] ), .COUT(
        \mult_23/CARRYB[13][1] ), .SUM(\mult_23/SUMB[13][1] ) );
  FADDER \mult_23/S1_13_0  ( .CIN(\mult_23/ab[13][0] ), .IN0(
        \mult_23/CARRYB[12][0] ), .IN1(\mult_23/SUMB[12][1] ), .COUT(
        \mult_23/CARRYB[13][0] ), .SUM(xy[13]) );
  FADDER \mult_23/S2_14_17  ( .CIN(\mult_23/ab[14][17] ), .IN0(
        \mult_23/CARRYB[13][17] ), .IN1(\mult_23/SUMB[13][18] ), .SUM(
        \mult_23/SUMB[14][17] ) );
  FADDER \mult_23/S2_14_16  ( .CIN(\mult_23/ab[14][16] ), .IN0(
        \mult_23/CARRYB[13][16] ), .IN1(\mult_23/SUMB[13][17] ), .COUT(
        \mult_23/CARRYB[14][16] ), .SUM(\mult_23/SUMB[14][16] ) );
  FADDER \mult_23/S2_14_15  ( .CIN(\mult_23/ab[14][15] ), .IN0(
        \mult_23/CARRYB[13][15] ), .IN1(\mult_23/SUMB[13][16] ), .COUT(
        \mult_23/CARRYB[14][15] ), .SUM(\mult_23/SUMB[14][15] ) );
  FADDER \mult_23/S2_14_14  ( .CIN(\mult_23/ab[14][14] ), .IN0(
        \mult_23/CARRYB[13][14] ), .IN1(\mult_23/SUMB[13][15] ), .COUT(
        \mult_23/CARRYB[14][14] ), .SUM(\mult_23/SUMB[14][14] ) );
  FADDER \mult_23/S2_14_13  ( .CIN(\mult_23/ab[14][13] ), .IN0(
        \mult_23/CARRYB[13][13] ), .IN1(\mult_23/SUMB[13][14] ), .COUT(
        \mult_23/CARRYB[14][13] ), .SUM(\mult_23/SUMB[14][13] ) );
  FADDER \mult_23/S2_14_12  ( .CIN(\mult_23/ab[14][12] ), .IN0(
        \mult_23/CARRYB[13][12] ), .IN1(\mult_23/SUMB[13][13] ), .COUT(
        \mult_23/CARRYB[14][12] ), .SUM(\mult_23/SUMB[14][12] ) );
  FADDER \mult_23/S2_14_11  ( .CIN(\mult_23/ab[14][11] ), .IN0(
        \mult_23/CARRYB[13][11] ), .IN1(\mult_23/SUMB[13][12] ), .COUT(
        \mult_23/CARRYB[14][11] ), .SUM(\mult_23/SUMB[14][11] ) );
  FADDER \mult_23/S2_14_10  ( .CIN(\mult_23/ab[14][10] ), .IN0(
        \mult_23/CARRYB[13][10] ), .IN1(\mult_23/SUMB[13][11] ), .COUT(
        \mult_23/CARRYB[14][10] ), .SUM(\mult_23/SUMB[14][10] ) );
  FADDER \mult_23/S2_14_9  ( .CIN(\mult_23/ab[14][9] ), .IN0(
        \mult_23/CARRYB[13][9] ), .IN1(\mult_23/SUMB[13][10] ), .COUT(
        \mult_23/CARRYB[14][9] ), .SUM(\mult_23/SUMB[14][9] ) );
  FADDER \mult_23/S2_14_8  ( .CIN(\mult_23/ab[14][8] ), .IN0(
        \mult_23/CARRYB[13][8] ), .IN1(\mult_23/SUMB[13][9] ), .COUT(
        \mult_23/CARRYB[14][8] ), .SUM(\mult_23/SUMB[14][8] ) );
  FADDER \mult_23/S2_14_7  ( .CIN(\mult_23/ab[14][7] ), .IN0(
        \mult_23/CARRYB[13][7] ), .IN1(\mult_23/SUMB[13][8] ), .COUT(
        \mult_23/CARRYB[14][7] ), .SUM(\mult_23/SUMB[14][7] ) );
  FADDER \mult_23/S2_14_6  ( .CIN(\mult_23/ab[14][6] ), .IN0(
        \mult_23/CARRYB[13][6] ), .IN1(\mult_23/SUMB[13][7] ), .COUT(
        \mult_23/CARRYB[14][6] ), .SUM(\mult_23/SUMB[14][6] ) );
  FADDER \mult_23/S2_14_5  ( .CIN(\mult_23/ab[14][5] ), .IN0(
        \mult_23/CARRYB[13][5] ), .IN1(\mult_23/SUMB[13][6] ), .COUT(
        \mult_23/CARRYB[14][5] ), .SUM(\mult_23/SUMB[14][5] ) );
  FADDER \mult_23/S2_14_4  ( .CIN(\mult_23/ab[14][4] ), .IN0(
        \mult_23/CARRYB[13][4] ), .IN1(\mult_23/SUMB[13][5] ), .COUT(
        \mult_23/CARRYB[14][4] ), .SUM(\mult_23/SUMB[14][4] ) );
  FADDER \mult_23/S2_14_3  ( .CIN(\mult_23/ab[14][3] ), .IN0(
        \mult_23/CARRYB[13][3] ), .IN1(\mult_23/SUMB[13][4] ), .COUT(
        \mult_23/CARRYB[14][3] ), .SUM(\mult_23/SUMB[14][3] ) );
  FADDER \mult_23/S2_14_2  ( .CIN(\mult_23/ab[14][2] ), .IN0(
        \mult_23/CARRYB[13][2] ), .IN1(\mult_23/SUMB[13][3] ), .COUT(
        \mult_23/CARRYB[14][2] ), .SUM(\mult_23/SUMB[14][2] ) );
  FADDER \mult_23/S2_14_1  ( .CIN(\mult_23/ab[14][1] ), .IN0(
        \mult_23/CARRYB[13][1] ), .IN1(\mult_23/SUMB[13][2] ), .COUT(
        \mult_23/CARRYB[14][1] ), .SUM(\mult_23/SUMB[14][1] ) );
  FADDER \mult_23/S1_14_0  ( .CIN(\mult_23/ab[14][0] ), .IN0(
        \mult_23/CARRYB[13][0] ), .IN1(\mult_23/SUMB[13][1] ), .COUT(
        \mult_23/CARRYB[14][0] ), .SUM(xy[14]) );
  FADDER \mult_23/S2_15_16  ( .CIN(\mult_23/ab[15][16] ), .IN0(
        \mult_23/CARRYB[14][16] ), .IN1(\mult_23/SUMB[14][17] ), .SUM(
        \mult_23/SUMB[15][16] ) );
  FADDER \mult_23/S2_15_15  ( .CIN(\mult_23/ab[15][15] ), .IN0(
        \mult_23/CARRYB[14][15] ), .IN1(\mult_23/SUMB[14][16] ), .COUT(
        \mult_23/CARRYB[15][15] ), .SUM(\mult_23/SUMB[15][15] ) );
  FADDER \mult_23/S2_15_14  ( .CIN(\mult_23/ab[15][14] ), .IN0(
        \mult_23/CARRYB[14][14] ), .IN1(\mult_23/SUMB[14][15] ), .COUT(
        \mult_23/CARRYB[15][14] ), .SUM(\mult_23/SUMB[15][14] ) );
  FADDER \mult_23/S2_15_13  ( .CIN(\mult_23/ab[15][13] ), .IN0(
        \mult_23/CARRYB[14][13] ), .IN1(\mult_23/SUMB[14][14] ), .COUT(
        \mult_23/CARRYB[15][13] ), .SUM(\mult_23/SUMB[15][13] ) );
  FADDER \mult_23/S2_15_12  ( .CIN(\mult_23/ab[15][12] ), .IN0(
        \mult_23/CARRYB[14][12] ), .IN1(\mult_23/SUMB[14][13] ), .COUT(
        \mult_23/CARRYB[15][12] ), .SUM(\mult_23/SUMB[15][12] ) );
  FADDER \mult_23/S2_15_11  ( .CIN(\mult_23/ab[15][11] ), .IN0(
        \mult_23/CARRYB[14][11] ), .IN1(\mult_23/SUMB[14][12] ), .COUT(
        \mult_23/CARRYB[15][11] ), .SUM(\mult_23/SUMB[15][11] ) );
  FADDER \mult_23/S2_15_10  ( .CIN(\mult_23/ab[15][10] ), .IN0(
        \mult_23/CARRYB[14][10] ), .IN1(\mult_23/SUMB[14][11] ), .COUT(
        \mult_23/CARRYB[15][10] ), .SUM(\mult_23/SUMB[15][10] ) );
  FADDER \mult_23/S2_15_9  ( .CIN(\mult_23/ab[15][9] ), .IN0(
        \mult_23/CARRYB[14][9] ), .IN1(\mult_23/SUMB[14][10] ), .COUT(
        \mult_23/CARRYB[15][9] ), .SUM(\mult_23/SUMB[15][9] ) );
  FADDER \mult_23/S2_15_8  ( .CIN(\mult_23/ab[15][8] ), .IN0(
        \mult_23/CARRYB[14][8] ), .IN1(\mult_23/SUMB[14][9] ), .COUT(
        \mult_23/CARRYB[15][8] ), .SUM(\mult_23/SUMB[15][8] ) );
  FADDER \mult_23/S2_15_7  ( .CIN(\mult_23/ab[15][7] ), .IN0(
        \mult_23/CARRYB[14][7] ), .IN1(\mult_23/SUMB[14][8] ), .COUT(
        \mult_23/CARRYB[15][7] ), .SUM(\mult_23/SUMB[15][7] ) );
  FADDER \mult_23/S2_15_6  ( .CIN(\mult_23/ab[15][6] ), .IN0(
        \mult_23/CARRYB[14][6] ), .IN1(\mult_23/SUMB[14][7] ), .COUT(
        \mult_23/CARRYB[15][6] ), .SUM(\mult_23/SUMB[15][6] ) );
  FADDER \mult_23/S2_15_5  ( .CIN(\mult_23/ab[15][5] ), .IN0(
        \mult_23/CARRYB[14][5] ), .IN1(\mult_23/SUMB[14][6] ), .COUT(
        \mult_23/CARRYB[15][5] ), .SUM(\mult_23/SUMB[15][5] ) );
  FADDER \mult_23/S2_15_4  ( .CIN(\mult_23/ab[15][4] ), .IN0(
        \mult_23/CARRYB[14][4] ), .IN1(\mult_23/SUMB[14][5] ), .COUT(
        \mult_23/CARRYB[15][4] ), .SUM(\mult_23/SUMB[15][4] ) );
  FADDER \mult_23/S2_15_3  ( .CIN(\mult_23/ab[15][3] ), .IN0(
        \mult_23/CARRYB[14][3] ), .IN1(\mult_23/SUMB[14][4] ), .COUT(
        \mult_23/CARRYB[15][3] ), .SUM(\mult_23/SUMB[15][3] ) );
  FADDER \mult_23/S2_15_2  ( .CIN(\mult_23/ab[15][2] ), .IN0(
        \mult_23/CARRYB[14][2] ), .IN1(\mult_23/SUMB[14][3] ), .COUT(
        \mult_23/CARRYB[15][2] ), .SUM(\mult_23/SUMB[15][2] ) );
  FADDER \mult_23/S2_15_1  ( .CIN(\mult_23/ab[15][1] ), .IN0(
        \mult_23/CARRYB[14][1] ), .IN1(\mult_23/SUMB[14][2] ), .COUT(
        \mult_23/CARRYB[15][1] ), .SUM(\mult_23/SUMB[15][1] ) );
  FADDER \mult_23/S1_15_0  ( .CIN(\mult_23/ab[15][0] ), .IN0(
        \mult_23/CARRYB[14][0] ), .IN1(\mult_23/SUMB[14][1] ), .COUT(
        \mult_23/CARRYB[15][0] ), .SUM(xy[15]) );
  FADDER \mult_23/S2_16_15  ( .CIN(\mult_23/ab[16][15] ), .IN0(
        \mult_23/CARRYB[15][15] ), .IN1(\mult_23/SUMB[15][16] ), .SUM(
        \mult_23/SUMB[16][15] ) );
  FADDER \mult_23/S2_16_14  ( .CIN(\mult_23/ab[16][14] ), .IN0(
        \mult_23/CARRYB[15][14] ), .IN1(\mult_23/SUMB[15][15] ), .COUT(
        \mult_23/CARRYB[16][14] ), .SUM(\mult_23/SUMB[16][14] ) );
  FADDER \mult_23/S2_16_13  ( .CIN(\mult_23/ab[16][13] ), .IN0(
        \mult_23/CARRYB[15][13] ), .IN1(\mult_23/SUMB[15][14] ), .COUT(
        \mult_23/CARRYB[16][13] ), .SUM(\mult_23/SUMB[16][13] ) );
  FADDER \mult_23/S2_16_12  ( .CIN(\mult_23/ab[16][12] ), .IN0(
        \mult_23/CARRYB[15][12] ), .IN1(\mult_23/SUMB[15][13] ), .COUT(
        \mult_23/CARRYB[16][12] ), .SUM(\mult_23/SUMB[16][12] ) );
  FADDER \mult_23/S2_16_11  ( .CIN(\mult_23/ab[16][11] ), .IN0(
        \mult_23/CARRYB[15][11] ), .IN1(\mult_23/SUMB[15][12] ), .COUT(
        \mult_23/CARRYB[16][11] ), .SUM(\mult_23/SUMB[16][11] ) );
  FADDER \mult_23/S2_16_10  ( .CIN(\mult_23/ab[16][10] ), .IN0(
        \mult_23/CARRYB[15][10] ), .IN1(\mult_23/SUMB[15][11] ), .COUT(
        \mult_23/CARRYB[16][10] ), .SUM(\mult_23/SUMB[16][10] ) );
  FADDER \mult_23/S2_16_9  ( .CIN(\mult_23/ab[16][9] ), .IN0(
        \mult_23/CARRYB[15][9] ), .IN1(\mult_23/SUMB[15][10] ), .COUT(
        \mult_23/CARRYB[16][9] ), .SUM(\mult_23/SUMB[16][9] ) );
  FADDER \mult_23/S2_16_8  ( .CIN(\mult_23/ab[16][8] ), .IN0(
        \mult_23/CARRYB[15][8] ), .IN1(\mult_23/SUMB[15][9] ), .COUT(
        \mult_23/CARRYB[16][8] ), .SUM(\mult_23/SUMB[16][8] ) );
  FADDER \mult_23/S2_16_7  ( .CIN(\mult_23/ab[16][7] ), .IN0(
        \mult_23/CARRYB[15][7] ), .IN1(\mult_23/SUMB[15][8] ), .COUT(
        \mult_23/CARRYB[16][7] ), .SUM(\mult_23/SUMB[16][7] ) );
  FADDER \mult_23/S2_16_6  ( .CIN(\mult_23/ab[16][6] ), .IN0(
        \mult_23/CARRYB[15][6] ), .IN1(\mult_23/SUMB[15][7] ), .COUT(
        \mult_23/CARRYB[16][6] ), .SUM(\mult_23/SUMB[16][6] ) );
  FADDER \mult_23/S2_16_5  ( .CIN(\mult_23/ab[16][5] ), .IN0(
        \mult_23/CARRYB[15][5] ), .IN1(\mult_23/SUMB[15][6] ), .COUT(
        \mult_23/CARRYB[16][5] ), .SUM(\mult_23/SUMB[16][5] ) );
  FADDER \mult_23/S2_16_4  ( .CIN(\mult_23/ab[16][4] ), .IN0(
        \mult_23/CARRYB[15][4] ), .IN1(\mult_23/SUMB[15][5] ), .COUT(
        \mult_23/CARRYB[16][4] ), .SUM(\mult_23/SUMB[16][4] ) );
  FADDER \mult_23/S2_16_3  ( .CIN(\mult_23/ab[16][3] ), .IN0(
        \mult_23/CARRYB[15][3] ), .IN1(\mult_23/SUMB[15][4] ), .COUT(
        \mult_23/CARRYB[16][3] ), .SUM(\mult_23/SUMB[16][3] ) );
  FADDER \mult_23/S2_16_2  ( .CIN(\mult_23/ab[16][2] ), .IN0(
        \mult_23/CARRYB[15][2] ), .IN1(\mult_23/SUMB[15][3] ), .COUT(
        \mult_23/CARRYB[16][2] ), .SUM(\mult_23/SUMB[16][2] ) );
  FADDER \mult_23/S2_16_1  ( .CIN(\mult_23/ab[16][1] ), .IN0(
        \mult_23/CARRYB[15][1] ), .IN1(\mult_23/SUMB[15][2] ), .COUT(
        \mult_23/CARRYB[16][1] ), .SUM(\mult_23/SUMB[16][1] ) );
  FADDER \mult_23/S1_16_0  ( .CIN(\mult_23/ab[16][0] ), .IN0(
        \mult_23/CARRYB[15][0] ), .IN1(\mult_23/SUMB[15][1] ), .COUT(
        \mult_23/CARRYB[16][0] ), .SUM(xy[16]) );
  FADDER \mult_23/S2_17_14  ( .CIN(\mult_23/ab[17][14] ), .IN0(
        \mult_23/CARRYB[16][14] ), .IN1(\mult_23/SUMB[16][15] ), .SUM(
        \mult_23/SUMB[17][14] ) );
  FADDER \mult_23/S2_17_13  ( .CIN(\mult_23/ab[17][13] ), .IN0(
        \mult_23/CARRYB[16][13] ), .IN1(\mult_23/SUMB[16][14] ), .COUT(
        \mult_23/CARRYB[17][13] ), .SUM(\mult_23/SUMB[17][13] ) );
  FADDER \mult_23/S2_17_12  ( .CIN(\mult_23/ab[17][12] ), .IN0(
        \mult_23/CARRYB[16][12] ), .IN1(\mult_23/SUMB[16][13] ), .COUT(
        \mult_23/CARRYB[17][12] ), .SUM(\mult_23/SUMB[17][12] ) );
  FADDER \mult_23/S2_17_11  ( .CIN(\mult_23/ab[17][11] ), .IN0(
        \mult_23/CARRYB[16][11] ), .IN1(\mult_23/SUMB[16][12] ), .COUT(
        \mult_23/CARRYB[17][11] ), .SUM(\mult_23/SUMB[17][11] ) );
  FADDER \mult_23/S2_17_10  ( .CIN(\mult_23/ab[17][10] ), .IN0(
        \mult_23/CARRYB[16][10] ), .IN1(\mult_23/SUMB[16][11] ), .COUT(
        \mult_23/CARRYB[17][10] ), .SUM(\mult_23/SUMB[17][10] ) );
  FADDER \mult_23/S2_17_9  ( .CIN(\mult_23/ab[17][9] ), .IN0(
        \mult_23/CARRYB[16][9] ), .IN1(\mult_23/SUMB[16][10] ), .COUT(
        \mult_23/CARRYB[17][9] ), .SUM(\mult_23/SUMB[17][9] ) );
  FADDER \mult_23/S2_17_8  ( .CIN(\mult_23/ab[17][8] ), .IN0(
        \mult_23/CARRYB[16][8] ), .IN1(\mult_23/SUMB[16][9] ), .COUT(
        \mult_23/CARRYB[17][8] ), .SUM(\mult_23/SUMB[17][8] ) );
  FADDER \mult_23/S2_17_7  ( .CIN(\mult_23/ab[17][7] ), .IN0(
        \mult_23/CARRYB[16][7] ), .IN1(\mult_23/SUMB[16][8] ), .COUT(
        \mult_23/CARRYB[17][7] ), .SUM(\mult_23/SUMB[17][7] ) );
  FADDER \mult_23/S2_17_6  ( .CIN(\mult_23/ab[17][6] ), .IN0(
        \mult_23/CARRYB[16][6] ), .IN1(\mult_23/SUMB[16][7] ), .COUT(
        \mult_23/CARRYB[17][6] ), .SUM(\mult_23/SUMB[17][6] ) );
  FADDER \mult_23/S2_17_5  ( .CIN(\mult_23/ab[17][5] ), .IN0(
        \mult_23/CARRYB[16][5] ), .IN1(\mult_23/SUMB[16][6] ), .COUT(
        \mult_23/CARRYB[17][5] ), .SUM(\mult_23/SUMB[17][5] ) );
  FADDER \mult_23/S2_17_4  ( .CIN(\mult_23/ab[17][4] ), .IN0(
        \mult_23/CARRYB[16][4] ), .IN1(\mult_23/SUMB[16][5] ), .COUT(
        \mult_23/CARRYB[17][4] ), .SUM(\mult_23/SUMB[17][4] ) );
  FADDER \mult_23/S2_17_3  ( .CIN(\mult_23/ab[17][3] ), .IN0(
        \mult_23/CARRYB[16][3] ), .IN1(\mult_23/SUMB[16][4] ), .COUT(
        \mult_23/CARRYB[17][3] ), .SUM(\mult_23/SUMB[17][3] ) );
  FADDER \mult_23/S2_17_2  ( .CIN(\mult_23/ab[17][2] ), .IN0(
        \mult_23/CARRYB[16][2] ), .IN1(\mult_23/SUMB[16][3] ), .COUT(
        \mult_23/CARRYB[17][2] ), .SUM(\mult_23/SUMB[17][2] ) );
  FADDER \mult_23/S2_17_1  ( .CIN(\mult_23/ab[17][1] ), .IN0(
        \mult_23/CARRYB[16][1] ), .IN1(\mult_23/SUMB[16][2] ), .COUT(
        \mult_23/CARRYB[17][1] ), .SUM(\mult_23/SUMB[17][1] ) );
  FADDER \mult_23/S1_17_0  ( .CIN(\mult_23/ab[17][0] ), .IN0(
        \mult_23/CARRYB[16][0] ), .IN1(\mult_23/SUMB[16][1] ), .COUT(
        \mult_23/CARRYB[17][0] ), .SUM(xy[17]) );
  FADDER \mult_23/S2_18_13  ( .CIN(\mult_23/ab[18][13] ), .IN0(
        \mult_23/CARRYB[17][13] ), .IN1(\mult_23/SUMB[17][14] ), .SUM(
        \mult_23/SUMB[18][13] ) );
  FADDER \mult_23/S2_18_12  ( .CIN(\mult_23/ab[18][12] ), .IN0(
        \mult_23/CARRYB[17][12] ), .IN1(\mult_23/SUMB[17][13] ), .COUT(
        \mult_23/CARRYB[18][12] ), .SUM(\mult_23/SUMB[18][12] ) );
  FADDER \mult_23/S2_18_11  ( .CIN(\mult_23/ab[18][11] ), .IN0(
        \mult_23/CARRYB[17][11] ), .IN1(\mult_23/SUMB[17][12] ), .COUT(
        \mult_23/CARRYB[18][11] ), .SUM(\mult_23/SUMB[18][11] ) );
  FADDER \mult_23/S2_18_10  ( .CIN(\mult_23/ab[18][10] ), .IN0(
        \mult_23/CARRYB[17][10] ), .IN1(\mult_23/SUMB[17][11] ), .COUT(
        \mult_23/CARRYB[18][10] ), .SUM(\mult_23/SUMB[18][10] ) );
  FADDER \mult_23/S2_18_9  ( .CIN(\mult_23/ab[18][9] ), .IN0(
        \mult_23/CARRYB[17][9] ), .IN1(\mult_23/SUMB[17][10] ), .COUT(
        \mult_23/CARRYB[18][9] ), .SUM(\mult_23/SUMB[18][9] ) );
  FADDER \mult_23/S2_18_8  ( .CIN(\mult_23/ab[18][8] ), .IN0(
        \mult_23/CARRYB[17][8] ), .IN1(\mult_23/SUMB[17][9] ), .COUT(
        \mult_23/CARRYB[18][8] ), .SUM(\mult_23/SUMB[18][8] ) );
  FADDER \mult_23/S2_18_7  ( .CIN(\mult_23/ab[18][7] ), .IN0(
        \mult_23/CARRYB[17][7] ), .IN1(\mult_23/SUMB[17][8] ), .COUT(
        \mult_23/CARRYB[18][7] ), .SUM(\mult_23/SUMB[18][7] ) );
  FADDER \mult_23/S2_18_6  ( .CIN(\mult_23/ab[18][6] ), .IN0(
        \mult_23/CARRYB[17][6] ), .IN1(\mult_23/SUMB[17][7] ), .COUT(
        \mult_23/CARRYB[18][6] ), .SUM(\mult_23/SUMB[18][6] ) );
  FADDER \mult_23/S2_18_5  ( .CIN(\mult_23/ab[18][5] ), .IN0(
        \mult_23/CARRYB[17][5] ), .IN1(\mult_23/SUMB[17][6] ), .COUT(
        \mult_23/CARRYB[18][5] ), .SUM(\mult_23/SUMB[18][5] ) );
  FADDER \mult_23/S2_18_4  ( .CIN(\mult_23/ab[18][4] ), .IN0(
        \mult_23/CARRYB[17][4] ), .IN1(\mult_23/SUMB[17][5] ), .COUT(
        \mult_23/CARRYB[18][4] ), .SUM(\mult_23/SUMB[18][4] ) );
  FADDER \mult_23/S2_18_3  ( .CIN(\mult_23/ab[18][3] ), .IN0(
        \mult_23/CARRYB[17][3] ), .IN1(\mult_23/SUMB[17][4] ), .COUT(
        \mult_23/CARRYB[18][3] ), .SUM(\mult_23/SUMB[18][3] ) );
  FADDER \mult_23/S2_18_2  ( .CIN(\mult_23/ab[18][2] ), .IN0(
        \mult_23/CARRYB[17][2] ), .IN1(\mult_23/SUMB[17][3] ), .COUT(
        \mult_23/CARRYB[18][2] ), .SUM(\mult_23/SUMB[18][2] ) );
  FADDER \mult_23/S2_18_1  ( .CIN(\mult_23/ab[18][1] ), .IN0(
        \mult_23/CARRYB[17][1] ), .IN1(\mult_23/SUMB[17][2] ), .COUT(
        \mult_23/CARRYB[18][1] ), .SUM(\mult_23/SUMB[18][1] ) );
  FADDER \mult_23/S1_18_0  ( .CIN(\mult_23/ab[18][0] ), .IN0(
        \mult_23/CARRYB[17][0] ), .IN1(\mult_23/SUMB[17][1] ), .COUT(
        \mult_23/CARRYB[18][0] ), .SUM(xy[18]) );
  FADDER \mult_23/S2_19_12  ( .CIN(\mult_23/ab[19][12] ), .IN0(
        \mult_23/CARRYB[18][12] ), .IN1(\mult_23/SUMB[18][13] ), .SUM(
        \mult_23/SUMB[19][12] ) );
  FADDER \mult_23/S2_19_11  ( .CIN(\mult_23/ab[19][11] ), .IN0(
        \mult_23/CARRYB[18][11] ), .IN1(\mult_23/SUMB[18][12] ), .COUT(
        \mult_23/CARRYB[19][11] ), .SUM(\mult_23/SUMB[19][11] ) );
  FADDER \mult_23/S2_19_10  ( .CIN(\mult_23/ab[19][10] ), .IN0(
        \mult_23/CARRYB[18][10] ), .IN1(\mult_23/SUMB[18][11] ), .COUT(
        \mult_23/CARRYB[19][10] ), .SUM(\mult_23/SUMB[19][10] ) );
  FADDER \mult_23/S2_19_9  ( .CIN(\mult_23/ab[19][9] ), .IN0(
        \mult_23/CARRYB[18][9] ), .IN1(\mult_23/SUMB[18][10] ), .COUT(
        \mult_23/CARRYB[19][9] ), .SUM(\mult_23/SUMB[19][9] ) );
  FADDER \mult_23/S2_19_8  ( .CIN(\mult_23/ab[19][8] ), .IN0(
        \mult_23/CARRYB[18][8] ), .IN1(\mult_23/SUMB[18][9] ), .COUT(
        \mult_23/CARRYB[19][8] ), .SUM(\mult_23/SUMB[19][8] ) );
  FADDER \mult_23/S2_19_7  ( .CIN(\mult_23/ab[19][7] ), .IN0(
        \mult_23/CARRYB[18][7] ), .IN1(\mult_23/SUMB[18][8] ), .COUT(
        \mult_23/CARRYB[19][7] ), .SUM(\mult_23/SUMB[19][7] ) );
  FADDER \mult_23/S2_19_6  ( .CIN(\mult_23/ab[19][6] ), .IN0(
        \mult_23/CARRYB[18][6] ), .IN1(\mult_23/SUMB[18][7] ), .COUT(
        \mult_23/CARRYB[19][6] ), .SUM(\mult_23/SUMB[19][6] ) );
  FADDER \mult_23/S2_19_5  ( .CIN(\mult_23/ab[19][5] ), .IN0(
        \mult_23/CARRYB[18][5] ), .IN1(\mult_23/SUMB[18][6] ), .COUT(
        \mult_23/CARRYB[19][5] ), .SUM(\mult_23/SUMB[19][5] ) );
  FADDER \mult_23/S2_19_4  ( .CIN(\mult_23/ab[19][4] ), .IN0(
        \mult_23/CARRYB[18][4] ), .IN1(\mult_23/SUMB[18][5] ), .COUT(
        \mult_23/CARRYB[19][4] ), .SUM(\mult_23/SUMB[19][4] ) );
  FADDER \mult_23/S2_19_3  ( .CIN(\mult_23/ab[19][3] ), .IN0(
        \mult_23/CARRYB[18][3] ), .IN1(\mult_23/SUMB[18][4] ), .COUT(
        \mult_23/CARRYB[19][3] ), .SUM(\mult_23/SUMB[19][3] ) );
  FADDER \mult_23/S2_19_2  ( .CIN(\mult_23/ab[19][2] ), .IN0(
        \mult_23/CARRYB[18][2] ), .IN1(\mult_23/SUMB[18][3] ), .COUT(
        \mult_23/CARRYB[19][2] ), .SUM(\mult_23/SUMB[19][2] ) );
  FADDER \mult_23/S2_19_1  ( .CIN(\mult_23/ab[19][1] ), .IN0(
        \mult_23/CARRYB[18][1] ), .IN1(\mult_23/SUMB[18][2] ), .COUT(
        \mult_23/CARRYB[19][1] ), .SUM(\mult_23/SUMB[19][1] ) );
  FADDER \mult_23/S1_19_0  ( .CIN(\mult_23/ab[19][0] ), .IN0(
        \mult_23/CARRYB[18][0] ), .IN1(\mult_23/SUMB[18][1] ), .COUT(
        \mult_23/CARRYB[19][0] ), .SUM(xy[19]) );
  FADDER \mult_23/S2_20_11  ( .CIN(\mult_23/ab[20][11] ), .IN0(
        \mult_23/CARRYB[19][11] ), .IN1(\mult_23/SUMB[19][12] ), .SUM(
        \mult_23/SUMB[20][11] ) );
  FADDER \mult_23/S2_20_10  ( .CIN(\mult_23/ab[20][10] ), .IN0(
        \mult_23/CARRYB[19][10] ), .IN1(\mult_23/SUMB[19][11] ), .COUT(
        \mult_23/CARRYB[20][10] ), .SUM(\mult_23/SUMB[20][10] ) );
  FADDER \mult_23/S2_20_9  ( .CIN(\mult_23/ab[20][9] ), .IN0(
        \mult_23/CARRYB[19][9] ), .IN1(\mult_23/SUMB[19][10] ), .COUT(
        \mult_23/CARRYB[20][9] ), .SUM(\mult_23/SUMB[20][9] ) );
  FADDER \mult_23/S2_20_8  ( .CIN(\mult_23/ab[20][8] ), .IN0(
        \mult_23/CARRYB[19][8] ), .IN1(\mult_23/SUMB[19][9] ), .COUT(
        \mult_23/CARRYB[20][8] ), .SUM(\mult_23/SUMB[20][8] ) );
  FADDER \mult_23/S2_20_7  ( .CIN(\mult_23/ab[20][7] ), .IN0(
        \mult_23/CARRYB[19][7] ), .IN1(\mult_23/SUMB[19][8] ), .COUT(
        \mult_23/CARRYB[20][7] ), .SUM(\mult_23/SUMB[20][7] ) );
  FADDER \mult_23/S2_20_6  ( .CIN(\mult_23/ab[20][6] ), .IN0(
        \mult_23/CARRYB[19][6] ), .IN1(\mult_23/SUMB[19][7] ), .COUT(
        \mult_23/CARRYB[20][6] ), .SUM(\mult_23/SUMB[20][6] ) );
  FADDER \mult_23/S2_20_5  ( .CIN(\mult_23/ab[20][5] ), .IN0(
        \mult_23/CARRYB[19][5] ), .IN1(\mult_23/SUMB[19][6] ), .COUT(
        \mult_23/CARRYB[20][5] ), .SUM(\mult_23/SUMB[20][5] ) );
  FADDER \mult_23/S2_20_4  ( .CIN(\mult_23/ab[20][4] ), .IN0(
        \mult_23/CARRYB[19][4] ), .IN1(\mult_23/SUMB[19][5] ), .COUT(
        \mult_23/CARRYB[20][4] ), .SUM(\mult_23/SUMB[20][4] ) );
  FADDER \mult_23/S2_20_3  ( .CIN(\mult_23/ab[20][3] ), .IN0(
        \mult_23/CARRYB[19][3] ), .IN1(\mult_23/SUMB[19][4] ), .COUT(
        \mult_23/CARRYB[20][3] ), .SUM(\mult_23/SUMB[20][3] ) );
  FADDER \mult_23/S2_20_2  ( .CIN(\mult_23/ab[20][2] ), .IN0(
        \mult_23/CARRYB[19][2] ), .IN1(\mult_23/SUMB[19][3] ), .COUT(
        \mult_23/CARRYB[20][2] ), .SUM(\mult_23/SUMB[20][2] ) );
  FADDER \mult_23/S2_20_1  ( .CIN(\mult_23/ab[20][1] ), .IN0(
        \mult_23/CARRYB[19][1] ), .IN1(\mult_23/SUMB[19][2] ), .COUT(
        \mult_23/CARRYB[20][1] ), .SUM(\mult_23/SUMB[20][1] ) );
  FADDER \mult_23/S1_20_0  ( .CIN(\mult_23/ab[20][0] ), .IN0(
        \mult_23/CARRYB[19][0] ), .IN1(\mult_23/SUMB[19][1] ), .COUT(
        \mult_23/CARRYB[20][0] ), .SUM(xy[20]) );
  FADDER \mult_23/S2_21_10  ( .CIN(\mult_23/ab[21][10] ), .IN0(
        \mult_23/CARRYB[20][10] ), .IN1(\mult_23/SUMB[20][11] ), .SUM(
        \mult_23/SUMB[21][10] ) );
  FADDER \mult_23/S2_21_9  ( .CIN(\mult_23/ab[21][9] ), .IN0(
        \mult_23/CARRYB[20][9] ), .IN1(\mult_23/SUMB[20][10] ), .COUT(
        \mult_23/CARRYB[21][9] ), .SUM(\mult_23/SUMB[21][9] ) );
  FADDER \mult_23/S2_21_8  ( .CIN(\mult_23/ab[21][8] ), .IN0(
        \mult_23/CARRYB[20][8] ), .IN1(\mult_23/SUMB[20][9] ), .COUT(
        \mult_23/CARRYB[21][8] ), .SUM(\mult_23/SUMB[21][8] ) );
  FADDER \mult_23/S2_21_7  ( .CIN(\mult_23/ab[21][7] ), .IN0(
        \mult_23/CARRYB[20][7] ), .IN1(\mult_23/SUMB[20][8] ), .COUT(
        \mult_23/CARRYB[21][7] ), .SUM(\mult_23/SUMB[21][7] ) );
  FADDER \mult_23/S2_21_6  ( .CIN(\mult_23/ab[21][6] ), .IN0(
        \mult_23/CARRYB[20][6] ), .IN1(\mult_23/SUMB[20][7] ), .COUT(
        \mult_23/CARRYB[21][6] ), .SUM(\mult_23/SUMB[21][6] ) );
  FADDER \mult_23/S2_21_5  ( .CIN(\mult_23/ab[21][5] ), .IN0(
        \mult_23/CARRYB[20][5] ), .IN1(\mult_23/SUMB[20][6] ), .COUT(
        \mult_23/CARRYB[21][5] ), .SUM(\mult_23/SUMB[21][5] ) );
  FADDER \mult_23/S2_21_4  ( .CIN(\mult_23/ab[21][4] ), .IN0(
        \mult_23/CARRYB[20][4] ), .IN1(\mult_23/SUMB[20][5] ), .COUT(
        \mult_23/CARRYB[21][4] ), .SUM(\mult_23/SUMB[21][4] ) );
  FADDER \mult_23/S2_21_3  ( .CIN(\mult_23/ab[21][3] ), .IN0(
        \mult_23/CARRYB[20][3] ), .IN1(\mult_23/SUMB[20][4] ), .COUT(
        \mult_23/CARRYB[21][3] ), .SUM(\mult_23/SUMB[21][3] ) );
  FADDER \mult_23/S2_21_2  ( .CIN(\mult_23/ab[21][2] ), .IN0(
        \mult_23/CARRYB[20][2] ), .IN1(\mult_23/SUMB[20][3] ), .COUT(
        \mult_23/CARRYB[21][2] ), .SUM(\mult_23/SUMB[21][2] ) );
  FADDER \mult_23/S2_21_1  ( .CIN(\mult_23/ab[21][1] ), .IN0(
        \mult_23/CARRYB[20][1] ), .IN1(\mult_23/SUMB[20][2] ), .COUT(
        \mult_23/CARRYB[21][1] ), .SUM(\mult_23/SUMB[21][1] ) );
  FADDER \mult_23/S1_21_0  ( .CIN(\mult_23/ab[21][0] ), .IN0(
        \mult_23/CARRYB[20][0] ), .IN1(\mult_23/SUMB[20][1] ), .COUT(
        \mult_23/CARRYB[21][0] ), .SUM(xy[21]) );
  FADDER \mult_23/S2_22_9  ( .CIN(\mult_23/ab[22][9] ), .IN0(
        \mult_23/CARRYB[21][9] ), .IN1(\mult_23/SUMB[21][10] ), .SUM(
        \mult_23/SUMB[22][9] ) );
  FADDER \mult_23/S2_22_8  ( .CIN(\mult_23/ab[22][8] ), .IN0(
        \mult_23/CARRYB[21][8] ), .IN1(\mult_23/SUMB[21][9] ), .COUT(
        \mult_23/CARRYB[22][8] ), .SUM(\mult_23/SUMB[22][8] ) );
  FADDER \mult_23/S2_22_7  ( .CIN(\mult_23/ab[22][7] ), .IN0(
        \mult_23/CARRYB[21][7] ), .IN1(\mult_23/SUMB[21][8] ), .COUT(
        \mult_23/CARRYB[22][7] ), .SUM(\mult_23/SUMB[22][7] ) );
  FADDER \mult_23/S2_22_6  ( .CIN(\mult_23/ab[22][6] ), .IN0(
        \mult_23/CARRYB[21][6] ), .IN1(\mult_23/SUMB[21][7] ), .COUT(
        \mult_23/CARRYB[22][6] ), .SUM(\mult_23/SUMB[22][6] ) );
  FADDER \mult_23/S2_22_5  ( .CIN(\mult_23/ab[22][5] ), .IN0(
        \mult_23/CARRYB[21][5] ), .IN1(\mult_23/SUMB[21][6] ), .COUT(
        \mult_23/CARRYB[22][5] ), .SUM(\mult_23/SUMB[22][5] ) );
  FADDER \mult_23/S2_22_4  ( .CIN(\mult_23/ab[22][4] ), .IN0(
        \mult_23/CARRYB[21][4] ), .IN1(\mult_23/SUMB[21][5] ), .COUT(
        \mult_23/CARRYB[22][4] ), .SUM(\mult_23/SUMB[22][4] ) );
  FADDER \mult_23/S2_22_3  ( .CIN(\mult_23/ab[22][3] ), .IN0(
        \mult_23/CARRYB[21][3] ), .IN1(\mult_23/SUMB[21][4] ), .COUT(
        \mult_23/CARRYB[22][3] ), .SUM(\mult_23/SUMB[22][3] ) );
  FADDER \mult_23/S2_22_2  ( .CIN(\mult_23/ab[22][2] ), .IN0(
        \mult_23/CARRYB[21][2] ), .IN1(\mult_23/SUMB[21][3] ), .COUT(
        \mult_23/CARRYB[22][2] ), .SUM(\mult_23/SUMB[22][2] ) );
  FADDER \mult_23/S2_22_1  ( .CIN(\mult_23/ab[22][1] ), .IN0(
        \mult_23/CARRYB[21][1] ), .IN1(\mult_23/SUMB[21][2] ), .COUT(
        \mult_23/CARRYB[22][1] ), .SUM(\mult_23/SUMB[22][1] ) );
  FADDER \mult_23/S1_22_0  ( .CIN(\mult_23/ab[22][0] ), .IN0(
        \mult_23/CARRYB[21][0] ), .IN1(\mult_23/SUMB[21][1] ), .COUT(
        \mult_23/CARRYB[22][0] ), .SUM(xy[22]) );
  FADDER \mult_23/S2_23_8  ( .CIN(\mult_23/ab[23][8] ), .IN0(
        \mult_23/CARRYB[22][8] ), .IN1(\mult_23/SUMB[22][9] ), .SUM(
        \mult_23/SUMB[23][8] ) );
  FADDER \mult_23/S2_23_7  ( .CIN(\mult_23/ab[23][7] ), .IN0(
        \mult_23/CARRYB[22][7] ), .IN1(\mult_23/SUMB[22][8] ), .COUT(
        \mult_23/CARRYB[23][7] ), .SUM(\mult_23/SUMB[23][7] ) );
  FADDER \mult_23/S2_23_6  ( .CIN(\mult_23/ab[23][6] ), .IN0(
        \mult_23/CARRYB[22][6] ), .IN1(\mult_23/SUMB[22][7] ), .COUT(
        \mult_23/CARRYB[23][6] ), .SUM(\mult_23/SUMB[23][6] ) );
  FADDER \mult_23/S2_23_5  ( .CIN(\mult_23/ab[23][5] ), .IN0(
        \mult_23/CARRYB[22][5] ), .IN1(\mult_23/SUMB[22][6] ), .COUT(
        \mult_23/CARRYB[23][5] ), .SUM(\mult_23/SUMB[23][5] ) );
  FADDER \mult_23/S2_23_4  ( .CIN(\mult_23/ab[23][4] ), .IN0(
        \mult_23/CARRYB[22][4] ), .IN1(\mult_23/SUMB[22][5] ), .COUT(
        \mult_23/CARRYB[23][4] ), .SUM(\mult_23/SUMB[23][4] ) );
  FADDER \mult_23/S2_23_3  ( .CIN(\mult_23/ab[23][3] ), .IN0(
        \mult_23/CARRYB[22][3] ), .IN1(\mult_23/SUMB[22][4] ), .COUT(
        \mult_23/CARRYB[23][3] ), .SUM(\mult_23/SUMB[23][3] ) );
  FADDER \mult_23/S2_23_2  ( .CIN(\mult_23/ab[23][2] ), .IN0(
        \mult_23/CARRYB[22][2] ), .IN1(\mult_23/SUMB[22][3] ), .COUT(
        \mult_23/CARRYB[23][2] ), .SUM(\mult_23/SUMB[23][2] ) );
  FADDER \mult_23/S2_23_1  ( .CIN(\mult_23/ab[23][1] ), .IN0(
        \mult_23/CARRYB[22][1] ), .IN1(\mult_23/SUMB[22][2] ), .COUT(
        \mult_23/CARRYB[23][1] ), .SUM(\mult_23/SUMB[23][1] ) );
  FADDER \mult_23/S1_23_0  ( .CIN(\mult_23/ab[23][0] ), .IN0(
        \mult_23/CARRYB[22][0] ), .IN1(\mult_23/SUMB[22][1] ), .COUT(
        \mult_23/CARRYB[23][0] ), .SUM(xy[23]) );
  FADDER \mult_23/S2_24_7  ( .CIN(\mult_23/ab[24][7] ), .IN0(
        \mult_23/CARRYB[23][7] ), .IN1(\mult_23/SUMB[23][8] ), .SUM(
        \mult_23/SUMB[24][7] ) );
  FADDER \mult_23/S2_24_6  ( .CIN(\mult_23/ab[24][6] ), .IN0(
        \mult_23/CARRYB[23][6] ), .IN1(\mult_23/SUMB[23][7] ), .COUT(
        \mult_23/CARRYB[24][6] ), .SUM(\mult_23/SUMB[24][6] ) );
  FADDER \mult_23/S2_24_5  ( .CIN(\mult_23/ab[24][5] ), .IN0(
        \mult_23/CARRYB[23][5] ), .IN1(\mult_23/SUMB[23][6] ), .COUT(
        \mult_23/CARRYB[24][5] ), .SUM(\mult_23/SUMB[24][5] ) );
  FADDER \mult_23/S2_24_4  ( .CIN(\mult_23/ab[24][4] ), .IN0(
        \mult_23/CARRYB[23][4] ), .IN1(\mult_23/SUMB[23][5] ), .COUT(
        \mult_23/CARRYB[24][4] ), .SUM(\mult_23/SUMB[24][4] ) );
  FADDER \mult_23/S2_24_3  ( .CIN(\mult_23/ab[24][3] ), .IN0(
        \mult_23/CARRYB[23][3] ), .IN1(\mult_23/SUMB[23][4] ), .COUT(
        \mult_23/CARRYB[24][3] ), .SUM(\mult_23/SUMB[24][3] ) );
  FADDER \mult_23/S2_24_2  ( .CIN(\mult_23/ab[24][2] ), .IN0(
        \mult_23/CARRYB[23][2] ), .IN1(\mult_23/SUMB[23][3] ), .COUT(
        \mult_23/CARRYB[24][2] ), .SUM(\mult_23/SUMB[24][2] ) );
  FADDER \mult_23/S2_24_1  ( .CIN(\mult_23/ab[24][1] ), .IN0(
        \mult_23/CARRYB[23][1] ), .IN1(\mult_23/SUMB[23][2] ), .COUT(
        \mult_23/CARRYB[24][1] ), .SUM(\mult_23/SUMB[24][1] ) );
  FADDER \mult_23/S1_24_0  ( .CIN(\mult_23/ab[24][0] ), .IN0(
        \mult_23/CARRYB[23][0] ), .IN1(\mult_23/SUMB[23][1] ), .COUT(
        \mult_23/CARRYB[24][0] ), .SUM(xy[24]) );
  FADDER \mult_23/S2_25_6  ( .CIN(\mult_23/ab[25][6] ), .IN0(
        \mult_23/CARRYB[24][6] ), .IN1(\mult_23/SUMB[24][7] ), .SUM(
        \mult_23/SUMB[25][6] ) );
  FADDER \mult_23/S2_25_5  ( .CIN(\mult_23/ab[25][5] ), .IN0(
        \mult_23/CARRYB[24][5] ), .IN1(\mult_23/SUMB[24][6] ), .COUT(
        \mult_23/CARRYB[25][5] ), .SUM(\mult_23/SUMB[25][5] ) );
  FADDER \mult_23/S2_25_4  ( .CIN(\mult_23/ab[25][4] ), .IN0(
        \mult_23/CARRYB[24][4] ), .IN1(\mult_23/SUMB[24][5] ), .COUT(
        \mult_23/CARRYB[25][4] ), .SUM(\mult_23/SUMB[25][4] ) );
  FADDER \mult_23/S2_25_3  ( .CIN(\mult_23/ab[25][3] ), .IN0(
        \mult_23/CARRYB[24][3] ), .IN1(\mult_23/SUMB[24][4] ), .COUT(
        \mult_23/CARRYB[25][3] ), .SUM(\mult_23/SUMB[25][3] ) );
  FADDER \mult_23/S2_25_2  ( .CIN(\mult_23/ab[25][2] ), .IN0(
        \mult_23/CARRYB[24][2] ), .IN1(\mult_23/SUMB[24][3] ), .COUT(
        \mult_23/CARRYB[25][2] ), .SUM(\mult_23/SUMB[25][2] ) );
  FADDER \mult_23/S2_25_1  ( .CIN(\mult_23/ab[25][1] ), .IN0(
        \mult_23/CARRYB[24][1] ), .IN1(\mult_23/SUMB[24][2] ), .COUT(
        \mult_23/CARRYB[25][1] ), .SUM(\mult_23/SUMB[25][1] ) );
  FADDER \mult_23/S1_25_0  ( .CIN(\mult_23/ab[25][0] ), .IN0(
        \mult_23/CARRYB[24][0] ), .IN1(\mult_23/SUMB[24][1] ), .COUT(
        \mult_23/CARRYB[25][0] ), .SUM(xy[25]) );
  FADDER \mult_23/S2_26_5  ( .CIN(\mult_23/ab[26][5] ), .IN0(
        \mult_23/CARRYB[25][5] ), .IN1(\mult_23/SUMB[25][6] ), .SUM(
        \mult_23/SUMB[26][5] ) );
  FADDER \mult_23/S2_26_4  ( .CIN(\mult_23/ab[26][4] ), .IN0(
        \mult_23/CARRYB[25][4] ), .IN1(\mult_23/SUMB[25][5] ), .COUT(
        \mult_23/CARRYB[26][4] ), .SUM(\mult_23/SUMB[26][4] ) );
  FADDER \mult_23/S2_26_3  ( .CIN(\mult_23/ab[26][3] ), .IN0(
        \mult_23/CARRYB[25][3] ), .IN1(\mult_23/SUMB[25][4] ), .COUT(
        \mult_23/CARRYB[26][3] ), .SUM(\mult_23/SUMB[26][3] ) );
  FADDER \mult_23/S2_26_2  ( .CIN(\mult_23/ab[26][2] ), .IN0(
        \mult_23/CARRYB[25][2] ), .IN1(\mult_23/SUMB[25][3] ), .COUT(
        \mult_23/CARRYB[26][2] ), .SUM(\mult_23/SUMB[26][2] ) );
  FADDER \mult_23/S2_26_1  ( .CIN(\mult_23/ab[26][1] ), .IN0(
        \mult_23/CARRYB[25][1] ), .IN1(\mult_23/SUMB[25][2] ), .COUT(
        \mult_23/CARRYB[26][1] ), .SUM(\mult_23/SUMB[26][1] ) );
  FADDER \mult_23/S1_26_0  ( .CIN(\mult_23/ab[26][0] ), .IN0(
        \mult_23/CARRYB[25][0] ), .IN1(\mult_23/SUMB[25][1] ), .COUT(
        \mult_23/CARRYB[26][0] ), .SUM(xy[26]) );
  FADDER \mult_23/S2_27_4  ( .CIN(\mult_23/ab[27][4] ), .IN0(
        \mult_23/CARRYB[26][4] ), .IN1(\mult_23/SUMB[26][5] ), .SUM(
        \mult_23/SUMB[27][4] ) );
  FADDER \mult_23/S2_27_3  ( .CIN(\mult_23/ab[27][3] ), .IN0(
        \mult_23/CARRYB[26][3] ), .IN1(\mult_23/SUMB[26][4] ), .COUT(
        \mult_23/CARRYB[27][3] ), .SUM(\mult_23/SUMB[27][3] ) );
  FADDER \mult_23/S2_27_2  ( .CIN(\mult_23/ab[27][2] ), .IN0(
        \mult_23/CARRYB[26][2] ), .IN1(\mult_23/SUMB[26][3] ), .COUT(
        \mult_23/CARRYB[27][2] ), .SUM(\mult_23/SUMB[27][2] ) );
  FADDER \mult_23/S2_27_1  ( .CIN(\mult_23/ab[27][1] ), .IN0(
        \mult_23/CARRYB[26][1] ), .IN1(\mult_23/SUMB[26][2] ), .COUT(
        \mult_23/CARRYB[27][1] ), .SUM(\mult_23/SUMB[27][1] ) );
  FADDER \mult_23/S1_27_0  ( .CIN(\mult_23/ab[27][0] ), .IN0(
        \mult_23/CARRYB[26][0] ), .IN1(\mult_23/SUMB[26][1] ), .COUT(
        \mult_23/CARRYB[27][0] ), .SUM(xy[27]) );
  FADDER \mult_23/S2_28_3  ( .CIN(\mult_23/ab[28][3] ), .IN0(
        \mult_23/CARRYB[27][3] ), .IN1(\mult_23/SUMB[27][4] ), .SUM(
        \mult_23/SUMB[28][3] ) );
  FADDER \mult_23/S2_28_2  ( .CIN(\mult_23/ab[28][2] ), .IN0(
        \mult_23/CARRYB[27][2] ), .IN1(\mult_23/SUMB[27][3] ), .COUT(
        \mult_23/CARRYB[28][2] ), .SUM(\mult_23/SUMB[28][2] ) );
  FADDER \mult_23/S2_28_1  ( .CIN(\mult_23/ab[28][1] ), .IN0(
        \mult_23/CARRYB[27][1] ), .IN1(\mult_23/SUMB[27][2] ), .COUT(
        \mult_23/CARRYB[28][1] ), .SUM(\mult_23/SUMB[28][1] ) );
  FADDER \mult_23/S1_28_0  ( .CIN(\mult_23/ab[28][0] ), .IN0(
        \mult_23/CARRYB[27][0] ), .IN1(\mult_23/SUMB[27][1] ), .COUT(
        \mult_23/CARRYB[28][0] ), .SUM(xy[28]) );
  FADDER \mult_23/S2_29_2  ( .CIN(\mult_23/ab[29][2] ), .IN0(
        \mult_23/CARRYB[28][2] ), .IN1(\mult_23/SUMB[28][3] ), .SUM(
        \mult_23/SUMB[29][2] ) );
  FADDER \mult_23/S2_29_1  ( .CIN(\mult_23/ab[29][1] ), .IN0(
        \mult_23/CARRYB[28][1] ), .IN1(\mult_23/SUMB[28][2] ), .COUT(
        \mult_23/CARRYB[29][1] ), .SUM(\mult_23/SUMB[29][1] ) );
  FADDER \mult_23/S1_29_0  ( .CIN(\mult_23/ab[29][0] ), .IN0(
        \mult_23/CARRYB[28][0] ), .IN1(\mult_23/SUMB[28][1] ), .COUT(
        \mult_23/CARRYB[29][0] ), .SUM(xy[29]) );
  FADDER \mult_23/S2_30_1  ( .CIN(\mult_23/ab[30][1] ), .IN0(
        \mult_23/CARRYB[29][1] ), .IN1(\mult_23/SUMB[29][2] ), .SUM(
        \mult_23/SUMB[30][1] ) );
  FADDER \mult_23/S1_30_0  ( .CIN(\mult_23/ab[30][0] ), .IN0(
        \mult_23/CARRYB[29][0] ), .IN1(\mult_23/SUMB[29][1] ), .COUT(
        \mult_23/CARRYB[30][0] ), .SUM(xy[30]) );
  FADDER \mult_23/S4_0  ( .CIN(\mult_23/ab[31][0] ), .IN0(
        \mult_23/CARRYB[30][0] ), .IN1(\mult_23/SUMB[30][1] ), .SUM(
        \mult_23/SUMB[31][0] ) );
  AND U37 ( .A(xy[0]), .B(o_reg[0]), .Z(\add_24/carry[1] ) );
  XOR U38 ( .A(o_reg[0]), .B(xy[0]), .Z(o[0]) );
  AND U39 ( .A(\mult_23/ab[0][1] ), .B(\mult_23/ab[1][0] ), .Z(
        \mult_23/CARRYB[1][0] ) );
  XOR U40 ( .A(\mult_23/ab[1][0] ), .B(\mult_23/ab[0][1] ), .Z(xy[1]) );
  AND U41 ( .A(\mult_23/ab[0][2] ), .B(\mult_23/ab[1][1] ), .Z(
        \mult_23/CARRYB[1][1] ) );
  XOR U42 ( .A(\mult_23/ab[1][1] ), .B(\mult_23/ab[0][2] ), .Z(
        \mult_23/SUMB[1][1] ) );
  AND U43 ( .A(\mult_23/ab[0][3] ), .B(\mult_23/ab[1][2] ), .Z(
        \mult_23/CARRYB[1][2] ) );
  XOR U44 ( .A(\mult_23/ab[1][2] ), .B(\mult_23/ab[0][3] ), .Z(
        \mult_23/SUMB[1][2] ) );
  AND U45 ( .A(\mult_23/ab[0][4] ), .B(\mult_23/ab[1][3] ), .Z(
        \mult_23/CARRYB[1][3] ) );
  XOR U46 ( .A(\mult_23/ab[1][3] ), .B(\mult_23/ab[0][4] ), .Z(
        \mult_23/SUMB[1][3] ) );
  AND U47 ( .A(\mult_23/ab[0][5] ), .B(\mult_23/ab[1][4] ), .Z(
        \mult_23/CARRYB[1][4] ) );
  XOR U48 ( .A(\mult_23/ab[1][4] ), .B(\mult_23/ab[0][5] ), .Z(
        \mult_23/SUMB[1][4] ) );
  AND U49 ( .A(\mult_23/ab[0][6] ), .B(\mult_23/ab[1][5] ), .Z(
        \mult_23/CARRYB[1][5] ) );
  XOR U50 ( .A(\mult_23/ab[1][5] ), .B(\mult_23/ab[0][6] ), .Z(
        \mult_23/SUMB[1][5] ) );
  AND U51 ( .A(\mult_23/ab[0][7] ), .B(\mult_23/ab[1][6] ), .Z(
        \mult_23/CARRYB[1][6] ) );
  XOR U52 ( .A(\mult_23/ab[1][6] ), .B(\mult_23/ab[0][7] ), .Z(
        \mult_23/SUMB[1][6] ) );
  AND U53 ( .A(\mult_23/ab[0][8] ), .B(\mult_23/ab[1][7] ), .Z(
        \mult_23/CARRYB[1][7] ) );
  XOR U54 ( .A(\mult_23/ab[1][7] ), .B(\mult_23/ab[0][8] ), .Z(
        \mult_23/SUMB[1][7] ) );
  AND U55 ( .A(\mult_23/ab[0][9] ), .B(\mult_23/ab[1][8] ), .Z(
        \mult_23/CARRYB[1][8] ) );
  XOR U56 ( .A(\mult_23/ab[1][8] ), .B(\mult_23/ab[0][9] ), .Z(
        \mult_23/SUMB[1][8] ) );
  AND U57 ( .A(\mult_23/ab[0][10] ), .B(\mult_23/ab[1][9] ), .Z(
        \mult_23/CARRYB[1][9] ) );
  XOR U58 ( .A(\mult_23/ab[1][9] ), .B(\mult_23/ab[0][10] ), .Z(
        \mult_23/SUMB[1][9] ) );
  AND U59 ( .A(\mult_23/ab[0][11] ), .B(\mult_23/ab[1][10] ), .Z(
        \mult_23/CARRYB[1][10] ) );
  XOR U60 ( .A(\mult_23/ab[1][10] ), .B(\mult_23/ab[0][11] ), .Z(
        \mult_23/SUMB[1][10] ) );
  AND U61 ( .A(\mult_23/ab[0][12] ), .B(\mult_23/ab[1][11] ), .Z(
        \mult_23/CARRYB[1][11] ) );
  XOR U62 ( .A(\mult_23/ab[1][11] ), .B(\mult_23/ab[0][12] ), .Z(
        \mult_23/SUMB[1][11] ) );
  AND U63 ( .A(\mult_23/ab[0][13] ), .B(\mult_23/ab[1][12] ), .Z(
        \mult_23/CARRYB[1][12] ) );
  XOR U64 ( .A(\mult_23/ab[1][12] ), .B(\mult_23/ab[0][13] ), .Z(
        \mult_23/SUMB[1][12] ) );
  AND U65 ( .A(\mult_23/ab[0][14] ), .B(\mult_23/ab[1][13] ), .Z(
        \mult_23/CARRYB[1][13] ) );
  XOR U66 ( .A(\mult_23/ab[1][13] ), .B(\mult_23/ab[0][14] ), .Z(
        \mult_23/SUMB[1][13] ) );
  AND U67 ( .A(\mult_23/ab[0][15] ), .B(\mult_23/ab[1][14] ), .Z(
        \mult_23/CARRYB[1][14] ) );
  XOR U68 ( .A(\mult_23/ab[1][14] ), .B(\mult_23/ab[0][15] ), .Z(
        \mult_23/SUMB[1][14] ) );
  AND U69 ( .A(\mult_23/ab[0][16] ), .B(\mult_23/ab[1][15] ), .Z(
        \mult_23/CARRYB[1][15] ) );
  XOR U70 ( .A(\mult_23/ab[1][15] ), .B(\mult_23/ab[0][16] ), .Z(
        \mult_23/SUMB[1][15] ) );
  AND U71 ( .A(\mult_23/ab[0][17] ), .B(\mult_23/ab[1][16] ), .Z(
        \mult_23/CARRYB[1][16] ) );
  XOR U72 ( .A(\mult_23/ab[1][16] ), .B(\mult_23/ab[0][17] ), .Z(
        \mult_23/SUMB[1][16] ) );
  AND U73 ( .A(\mult_23/ab[0][18] ), .B(\mult_23/ab[1][17] ), .Z(
        \mult_23/CARRYB[1][17] ) );
  XOR U74 ( .A(\mult_23/ab[1][17] ), .B(\mult_23/ab[0][18] ), .Z(
        \mult_23/SUMB[1][17] ) );
  AND U75 ( .A(\mult_23/ab[0][19] ), .B(\mult_23/ab[1][18] ), .Z(
        \mult_23/CARRYB[1][18] ) );
  XOR U76 ( .A(\mult_23/ab[1][18] ), .B(\mult_23/ab[0][19] ), .Z(
        \mult_23/SUMB[1][18] ) );
  AND U77 ( .A(\mult_23/ab[0][20] ), .B(\mult_23/ab[1][19] ), .Z(
        \mult_23/CARRYB[1][19] ) );
  XOR U78 ( .A(\mult_23/ab[1][19] ), .B(\mult_23/ab[0][20] ), .Z(
        \mult_23/SUMB[1][19] ) );
  AND U79 ( .A(\mult_23/ab[0][21] ), .B(\mult_23/ab[1][20] ), .Z(
        \mult_23/CARRYB[1][20] ) );
  XOR U80 ( .A(\mult_23/ab[1][20] ), .B(\mult_23/ab[0][21] ), .Z(
        \mult_23/SUMB[1][20] ) );
  AND U81 ( .A(\mult_23/ab[0][22] ), .B(\mult_23/ab[1][21] ), .Z(
        \mult_23/CARRYB[1][21] ) );
  XOR U82 ( .A(\mult_23/ab[1][21] ), .B(\mult_23/ab[0][22] ), .Z(
        \mult_23/SUMB[1][21] ) );
  AND U83 ( .A(\mult_23/ab[0][23] ), .B(\mult_23/ab[1][22] ), .Z(
        \mult_23/CARRYB[1][22] ) );
  XOR U84 ( .A(\mult_23/ab[1][22] ), .B(\mult_23/ab[0][23] ), .Z(
        \mult_23/SUMB[1][22] ) );
  AND U85 ( .A(\mult_23/ab[0][24] ), .B(\mult_23/ab[1][23] ), .Z(
        \mult_23/CARRYB[1][23] ) );
  XOR U86 ( .A(\mult_23/ab[1][23] ), .B(\mult_23/ab[0][24] ), .Z(
        \mult_23/SUMB[1][23] ) );
  AND U87 ( .A(\mult_23/ab[0][25] ), .B(\mult_23/ab[1][24] ), .Z(
        \mult_23/CARRYB[1][24] ) );
  XOR U88 ( .A(\mult_23/ab[1][24] ), .B(\mult_23/ab[0][25] ), .Z(
        \mult_23/SUMB[1][24] ) );
  AND U89 ( .A(\mult_23/ab[0][26] ), .B(\mult_23/ab[1][25] ), .Z(
        \mult_23/CARRYB[1][25] ) );
  XOR U90 ( .A(\mult_23/ab[1][25] ), .B(\mult_23/ab[0][26] ), .Z(
        \mult_23/SUMB[1][25] ) );
  AND U91 ( .A(\mult_23/ab[0][27] ), .B(\mult_23/ab[1][26] ), .Z(
        \mult_23/CARRYB[1][26] ) );
  XOR U92 ( .A(\mult_23/ab[1][26] ), .B(\mult_23/ab[0][27] ), .Z(
        \mult_23/SUMB[1][26] ) );
  AND U93 ( .A(\mult_23/ab[0][28] ), .B(\mult_23/ab[1][27] ), .Z(
        \mult_23/CARRYB[1][27] ) );
  XOR U94 ( .A(\mult_23/ab[1][27] ), .B(\mult_23/ab[0][28] ), .Z(
        \mult_23/SUMB[1][27] ) );
  AND U95 ( .A(\mult_23/ab[0][29] ), .B(\mult_23/ab[1][28] ), .Z(
        \mult_23/CARRYB[1][28] ) );
  XOR U96 ( .A(\mult_23/ab[1][28] ), .B(\mult_23/ab[0][29] ), .Z(
        \mult_23/SUMB[1][28] ) );
  AND U97 ( .A(\mult_23/ab[0][30] ), .B(\mult_23/ab[1][29] ), .Z(
        \mult_23/CARRYB[1][29] ) );
  XOR U98 ( .A(\mult_23/ab[1][29] ), .B(\mult_23/ab[0][30] ), .Z(
        \mult_23/SUMB[1][29] ) );
  XOR U99 ( .A(\mult_23/ab[0][31] ), .B(\mult_23/ab[1][30] ), .Z(
        \mult_23/SUMB[1][30] ) );
  AND U100 ( .A(e_input[0]), .B(g_input[0]), .Z(xy[0]) );
  AND U101 ( .A(e_input[9]), .B(g_input[9]), .Z(\mult_23/ab[9][9] ) );
  AND U102 ( .A(g_input[9]), .B(e_input[8]), .Z(\mult_23/ab[9][8] ) );
  AND U103 ( .A(g_input[9]), .B(e_input[7]), .Z(\mult_23/ab[9][7] ) );
  AND U104 ( .A(g_input[9]), .B(e_input[6]), .Z(\mult_23/ab[9][6] ) );
  AND U105 ( .A(g_input[9]), .B(e_input[5]), .Z(\mult_23/ab[9][5] ) );
  AND U106 ( .A(g_input[9]), .B(e_input[4]), .Z(\mult_23/ab[9][4] ) );
  AND U107 ( .A(g_input[9]), .B(e_input[3]), .Z(\mult_23/ab[9][3] ) );
  AND U108 ( .A(g_input[9]), .B(e_input[2]), .Z(\mult_23/ab[9][2] ) );
  AND U109 ( .A(g_input[9]), .B(e_input[22]), .Z(\mult_23/ab[9][22] ) );
  AND U110 ( .A(g_input[9]), .B(e_input[21]), .Z(\mult_23/ab[9][21] ) );
  AND U111 ( .A(g_input[9]), .B(e_input[20]), .Z(\mult_23/ab[9][20] ) );
  AND U112 ( .A(g_input[9]), .B(e_input[1]), .Z(\mult_23/ab[9][1] ) );
  AND U113 ( .A(g_input[9]), .B(e_input[19]), .Z(\mult_23/ab[9][19] ) );
  AND U114 ( .A(g_input[9]), .B(e_input[18]), .Z(\mult_23/ab[9][18] ) );
  AND U115 ( .A(g_input[9]), .B(e_input[17]), .Z(\mult_23/ab[9][17] ) );
  AND U116 ( .A(g_input[9]), .B(e_input[16]), .Z(\mult_23/ab[9][16] ) );
  AND U117 ( .A(g_input[9]), .B(e_input[15]), .Z(\mult_23/ab[9][15] ) );
  AND U118 ( .A(g_input[9]), .B(e_input[14]), .Z(\mult_23/ab[9][14] ) );
  AND U119 ( .A(g_input[9]), .B(e_input[13]), .Z(\mult_23/ab[9][13] ) );
  AND U120 ( .A(g_input[9]), .B(e_input[12]), .Z(\mult_23/ab[9][12] ) );
  AND U121 ( .A(g_input[9]), .B(e_input[11]), .Z(\mult_23/ab[9][11] ) );
  AND U122 ( .A(g_input[9]), .B(e_input[10]), .Z(\mult_23/ab[9][10] ) );
  AND U123 ( .A(e_input[0]), .B(g_input[9]), .Z(\mult_23/ab[9][0] ) );
  AND U124 ( .A(e_input[9]), .B(g_input[8]), .Z(\mult_23/ab[8][9] ) );
  AND U125 ( .A(e_input[8]), .B(g_input[8]), .Z(\mult_23/ab[8][8] ) );
  AND U126 ( .A(e_input[7]), .B(g_input[8]), .Z(\mult_23/ab[8][7] ) );
  AND U127 ( .A(e_input[6]), .B(g_input[8]), .Z(\mult_23/ab[8][6] ) );
  AND U128 ( .A(e_input[5]), .B(g_input[8]), .Z(\mult_23/ab[8][5] ) );
  AND U129 ( .A(e_input[4]), .B(g_input[8]), .Z(\mult_23/ab[8][4] ) );
  AND U130 ( .A(e_input[3]), .B(g_input[8]), .Z(\mult_23/ab[8][3] ) );
  AND U131 ( .A(e_input[2]), .B(g_input[8]), .Z(\mult_23/ab[8][2] ) );
  AND U132 ( .A(g_input[8]), .B(e_input[23]), .Z(\mult_23/ab[8][23] ) );
  AND U133 ( .A(e_input[22]), .B(g_input[8]), .Z(\mult_23/ab[8][22] ) );
  AND U134 ( .A(e_input[21]), .B(g_input[8]), .Z(\mult_23/ab[8][21] ) );
  AND U135 ( .A(e_input[20]), .B(g_input[8]), .Z(\mult_23/ab[8][20] ) );
  AND U136 ( .A(e_input[1]), .B(g_input[8]), .Z(\mult_23/ab[8][1] ) );
  AND U137 ( .A(e_input[19]), .B(g_input[8]), .Z(\mult_23/ab[8][19] ) );
  AND U138 ( .A(e_input[18]), .B(g_input[8]), .Z(\mult_23/ab[8][18] ) );
  AND U139 ( .A(e_input[17]), .B(g_input[8]), .Z(\mult_23/ab[8][17] ) );
  AND U140 ( .A(e_input[16]), .B(g_input[8]), .Z(\mult_23/ab[8][16] ) );
  AND U141 ( .A(e_input[15]), .B(g_input[8]), .Z(\mult_23/ab[8][15] ) );
  AND U142 ( .A(e_input[14]), .B(g_input[8]), .Z(\mult_23/ab[8][14] ) );
  AND U143 ( .A(e_input[13]), .B(g_input[8]), .Z(\mult_23/ab[8][13] ) );
  AND U144 ( .A(e_input[12]), .B(g_input[8]), .Z(\mult_23/ab[8][12] ) );
  AND U145 ( .A(e_input[11]), .B(g_input[8]), .Z(\mult_23/ab[8][11] ) );
  AND U146 ( .A(e_input[10]), .B(g_input[8]), .Z(\mult_23/ab[8][10] ) );
  AND U147 ( .A(e_input[0]), .B(g_input[8]), .Z(\mult_23/ab[8][0] ) );
  AND U148 ( .A(e_input[9]), .B(g_input[7]), .Z(\mult_23/ab[7][9] ) );
  AND U149 ( .A(e_input[8]), .B(g_input[7]), .Z(\mult_23/ab[7][8] ) );
  AND U150 ( .A(e_input[7]), .B(g_input[7]), .Z(\mult_23/ab[7][7] ) );
  AND U151 ( .A(e_input[6]), .B(g_input[7]), .Z(\mult_23/ab[7][6] ) );
  AND U152 ( .A(e_input[5]), .B(g_input[7]), .Z(\mult_23/ab[7][5] ) );
  AND U153 ( .A(e_input[4]), .B(g_input[7]), .Z(\mult_23/ab[7][4] ) );
  AND U154 ( .A(e_input[3]), .B(g_input[7]), .Z(\mult_23/ab[7][3] ) );
  AND U155 ( .A(e_input[2]), .B(g_input[7]), .Z(\mult_23/ab[7][2] ) );
  AND U156 ( .A(g_input[7]), .B(e_input[24]), .Z(\mult_23/ab[7][24] ) );
  AND U157 ( .A(e_input[23]), .B(g_input[7]), .Z(\mult_23/ab[7][23] ) );
  AND U158 ( .A(e_input[22]), .B(g_input[7]), .Z(\mult_23/ab[7][22] ) );
  AND U159 ( .A(e_input[21]), .B(g_input[7]), .Z(\mult_23/ab[7][21] ) );
  AND U160 ( .A(e_input[20]), .B(g_input[7]), .Z(\mult_23/ab[7][20] ) );
  AND U161 ( .A(e_input[1]), .B(g_input[7]), .Z(\mult_23/ab[7][1] ) );
  AND U162 ( .A(e_input[19]), .B(g_input[7]), .Z(\mult_23/ab[7][19] ) );
  AND U163 ( .A(e_input[18]), .B(g_input[7]), .Z(\mult_23/ab[7][18] ) );
  AND U164 ( .A(e_input[17]), .B(g_input[7]), .Z(\mult_23/ab[7][17] ) );
  AND U165 ( .A(e_input[16]), .B(g_input[7]), .Z(\mult_23/ab[7][16] ) );
  AND U166 ( .A(e_input[15]), .B(g_input[7]), .Z(\mult_23/ab[7][15] ) );
  AND U167 ( .A(e_input[14]), .B(g_input[7]), .Z(\mult_23/ab[7][14] ) );
  AND U168 ( .A(e_input[13]), .B(g_input[7]), .Z(\mult_23/ab[7][13] ) );
  AND U169 ( .A(e_input[12]), .B(g_input[7]), .Z(\mult_23/ab[7][12] ) );
  AND U170 ( .A(e_input[11]), .B(g_input[7]), .Z(\mult_23/ab[7][11] ) );
  AND U171 ( .A(e_input[10]), .B(g_input[7]), .Z(\mult_23/ab[7][10] ) );
  AND U172 ( .A(e_input[0]), .B(g_input[7]), .Z(\mult_23/ab[7][0] ) );
  AND U173 ( .A(e_input[9]), .B(g_input[6]), .Z(\mult_23/ab[6][9] ) );
  AND U174 ( .A(e_input[8]), .B(g_input[6]), .Z(\mult_23/ab[6][8] ) );
  AND U175 ( .A(e_input[7]), .B(g_input[6]), .Z(\mult_23/ab[6][7] ) );
  AND U176 ( .A(e_input[6]), .B(g_input[6]), .Z(\mult_23/ab[6][6] ) );
  AND U177 ( .A(e_input[5]), .B(g_input[6]), .Z(\mult_23/ab[6][5] ) );
  AND U178 ( .A(e_input[4]), .B(g_input[6]), .Z(\mult_23/ab[6][4] ) );
  AND U179 ( .A(e_input[3]), .B(g_input[6]), .Z(\mult_23/ab[6][3] ) );
  AND U180 ( .A(e_input[2]), .B(g_input[6]), .Z(\mult_23/ab[6][2] ) );
  AND U181 ( .A(g_input[6]), .B(e_input[25]), .Z(\mult_23/ab[6][25] ) );
  AND U182 ( .A(e_input[24]), .B(g_input[6]), .Z(\mult_23/ab[6][24] ) );
  AND U183 ( .A(e_input[23]), .B(g_input[6]), .Z(\mult_23/ab[6][23] ) );
  AND U184 ( .A(e_input[22]), .B(g_input[6]), .Z(\mult_23/ab[6][22] ) );
  AND U185 ( .A(e_input[21]), .B(g_input[6]), .Z(\mult_23/ab[6][21] ) );
  AND U186 ( .A(e_input[20]), .B(g_input[6]), .Z(\mult_23/ab[6][20] ) );
  AND U187 ( .A(e_input[1]), .B(g_input[6]), .Z(\mult_23/ab[6][1] ) );
  AND U188 ( .A(e_input[19]), .B(g_input[6]), .Z(\mult_23/ab[6][19] ) );
  AND U189 ( .A(e_input[18]), .B(g_input[6]), .Z(\mult_23/ab[6][18] ) );
  AND U190 ( .A(e_input[17]), .B(g_input[6]), .Z(\mult_23/ab[6][17] ) );
  AND U191 ( .A(e_input[16]), .B(g_input[6]), .Z(\mult_23/ab[6][16] ) );
  AND U192 ( .A(e_input[15]), .B(g_input[6]), .Z(\mult_23/ab[6][15] ) );
  AND U193 ( .A(e_input[14]), .B(g_input[6]), .Z(\mult_23/ab[6][14] ) );
  AND U194 ( .A(e_input[13]), .B(g_input[6]), .Z(\mult_23/ab[6][13] ) );
  AND U195 ( .A(e_input[12]), .B(g_input[6]), .Z(\mult_23/ab[6][12] ) );
  AND U196 ( .A(e_input[11]), .B(g_input[6]), .Z(\mult_23/ab[6][11] ) );
  AND U197 ( .A(e_input[10]), .B(g_input[6]), .Z(\mult_23/ab[6][10] ) );
  AND U198 ( .A(e_input[0]), .B(g_input[6]), .Z(\mult_23/ab[6][0] ) );
  AND U199 ( .A(e_input[9]), .B(g_input[5]), .Z(\mult_23/ab[5][9] ) );
  AND U200 ( .A(e_input[8]), .B(g_input[5]), .Z(\mult_23/ab[5][8] ) );
  AND U201 ( .A(e_input[7]), .B(g_input[5]), .Z(\mult_23/ab[5][7] ) );
  AND U202 ( .A(e_input[6]), .B(g_input[5]), .Z(\mult_23/ab[5][6] ) );
  AND U203 ( .A(e_input[5]), .B(g_input[5]), .Z(\mult_23/ab[5][5] ) );
  AND U204 ( .A(e_input[4]), .B(g_input[5]), .Z(\mult_23/ab[5][4] ) );
  AND U205 ( .A(e_input[3]), .B(g_input[5]), .Z(\mult_23/ab[5][3] ) );
  AND U206 ( .A(e_input[2]), .B(g_input[5]), .Z(\mult_23/ab[5][2] ) );
  AND U207 ( .A(g_input[5]), .B(e_input[26]), .Z(\mult_23/ab[5][26] ) );
  AND U208 ( .A(e_input[25]), .B(g_input[5]), .Z(\mult_23/ab[5][25] ) );
  AND U209 ( .A(e_input[24]), .B(g_input[5]), .Z(\mult_23/ab[5][24] ) );
  AND U210 ( .A(e_input[23]), .B(g_input[5]), .Z(\mult_23/ab[5][23] ) );
  AND U211 ( .A(e_input[22]), .B(g_input[5]), .Z(\mult_23/ab[5][22] ) );
  AND U212 ( .A(e_input[21]), .B(g_input[5]), .Z(\mult_23/ab[5][21] ) );
  AND U213 ( .A(e_input[20]), .B(g_input[5]), .Z(\mult_23/ab[5][20] ) );
  AND U214 ( .A(e_input[1]), .B(g_input[5]), .Z(\mult_23/ab[5][1] ) );
  AND U215 ( .A(e_input[19]), .B(g_input[5]), .Z(\mult_23/ab[5][19] ) );
  AND U216 ( .A(e_input[18]), .B(g_input[5]), .Z(\mult_23/ab[5][18] ) );
  AND U217 ( .A(e_input[17]), .B(g_input[5]), .Z(\mult_23/ab[5][17] ) );
  AND U218 ( .A(e_input[16]), .B(g_input[5]), .Z(\mult_23/ab[5][16] ) );
  AND U219 ( .A(e_input[15]), .B(g_input[5]), .Z(\mult_23/ab[5][15] ) );
  AND U220 ( .A(e_input[14]), .B(g_input[5]), .Z(\mult_23/ab[5][14] ) );
  AND U221 ( .A(e_input[13]), .B(g_input[5]), .Z(\mult_23/ab[5][13] ) );
  AND U222 ( .A(e_input[12]), .B(g_input[5]), .Z(\mult_23/ab[5][12] ) );
  AND U223 ( .A(e_input[11]), .B(g_input[5]), .Z(\mult_23/ab[5][11] ) );
  AND U224 ( .A(e_input[10]), .B(g_input[5]), .Z(\mult_23/ab[5][10] ) );
  AND U225 ( .A(e_input[0]), .B(g_input[5]), .Z(\mult_23/ab[5][0] ) );
  AND U226 ( .A(e_input[9]), .B(g_input[4]), .Z(\mult_23/ab[4][9] ) );
  AND U227 ( .A(e_input[8]), .B(g_input[4]), .Z(\mult_23/ab[4][8] ) );
  AND U228 ( .A(e_input[7]), .B(g_input[4]), .Z(\mult_23/ab[4][7] ) );
  AND U229 ( .A(e_input[6]), .B(g_input[4]), .Z(\mult_23/ab[4][6] ) );
  AND U230 ( .A(e_input[5]), .B(g_input[4]), .Z(\mult_23/ab[4][5] ) );
  AND U231 ( .A(e_input[4]), .B(g_input[4]), .Z(\mult_23/ab[4][4] ) );
  AND U232 ( .A(e_input[3]), .B(g_input[4]), .Z(\mult_23/ab[4][3] ) );
  AND U233 ( .A(e_input[2]), .B(g_input[4]), .Z(\mult_23/ab[4][2] ) );
  AND U234 ( .A(g_input[4]), .B(e_input[27]), .Z(\mult_23/ab[4][27] ) );
  AND U235 ( .A(e_input[26]), .B(g_input[4]), .Z(\mult_23/ab[4][26] ) );
  AND U236 ( .A(e_input[25]), .B(g_input[4]), .Z(\mult_23/ab[4][25] ) );
  AND U237 ( .A(e_input[24]), .B(g_input[4]), .Z(\mult_23/ab[4][24] ) );
  AND U238 ( .A(e_input[23]), .B(g_input[4]), .Z(\mult_23/ab[4][23] ) );
  AND U239 ( .A(e_input[22]), .B(g_input[4]), .Z(\mult_23/ab[4][22] ) );
  AND U240 ( .A(e_input[21]), .B(g_input[4]), .Z(\mult_23/ab[4][21] ) );
  AND U241 ( .A(e_input[20]), .B(g_input[4]), .Z(\mult_23/ab[4][20] ) );
  AND U242 ( .A(e_input[1]), .B(g_input[4]), .Z(\mult_23/ab[4][1] ) );
  AND U243 ( .A(e_input[19]), .B(g_input[4]), .Z(\mult_23/ab[4][19] ) );
  AND U244 ( .A(e_input[18]), .B(g_input[4]), .Z(\mult_23/ab[4][18] ) );
  AND U245 ( .A(e_input[17]), .B(g_input[4]), .Z(\mult_23/ab[4][17] ) );
  AND U246 ( .A(e_input[16]), .B(g_input[4]), .Z(\mult_23/ab[4][16] ) );
  AND U247 ( .A(e_input[15]), .B(g_input[4]), .Z(\mult_23/ab[4][15] ) );
  AND U248 ( .A(e_input[14]), .B(g_input[4]), .Z(\mult_23/ab[4][14] ) );
  AND U249 ( .A(e_input[13]), .B(g_input[4]), .Z(\mult_23/ab[4][13] ) );
  AND U250 ( .A(e_input[12]), .B(g_input[4]), .Z(\mult_23/ab[4][12] ) );
  AND U251 ( .A(e_input[11]), .B(g_input[4]), .Z(\mult_23/ab[4][11] ) );
  AND U252 ( .A(e_input[10]), .B(g_input[4]), .Z(\mult_23/ab[4][10] ) );
  AND U253 ( .A(e_input[0]), .B(g_input[4]), .Z(\mult_23/ab[4][0] ) );
  AND U254 ( .A(e_input[9]), .B(g_input[3]), .Z(\mult_23/ab[3][9] ) );
  AND U255 ( .A(e_input[8]), .B(g_input[3]), .Z(\mult_23/ab[3][8] ) );
  AND U256 ( .A(e_input[7]), .B(g_input[3]), .Z(\mult_23/ab[3][7] ) );
  AND U257 ( .A(e_input[6]), .B(g_input[3]), .Z(\mult_23/ab[3][6] ) );
  AND U258 ( .A(e_input[5]), .B(g_input[3]), .Z(\mult_23/ab[3][5] ) );
  AND U259 ( .A(e_input[4]), .B(g_input[3]), .Z(\mult_23/ab[3][4] ) );
  AND U260 ( .A(e_input[3]), .B(g_input[3]), .Z(\mult_23/ab[3][3] ) );
  AND U261 ( .A(e_input[2]), .B(g_input[3]), .Z(\mult_23/ab[3][2] ) );
  AND U262 ( .A(g_input[3]), .B(e_input[28]), .Z(\mult_23/ab[3][28] ) );
  AND U263 ( .A(e_input[27]), .B(g_input[3]), .Z(\mult_23/ab[3][27] ) );
  AND U264 ( .A(e_input[26]), .B(g_input[3]), .Z(\mult_23/ab[3][26] ) );
  AND U265 ( .A(e_input[25]), .B(g_input[3]), .Z(\mult_23/ab[3][25] ) );
  AND U266 ( .A(e_input[24]), .B(g_input[3]), .Z(\mult_23/ab[3][24] ) );
  AND U267 ( .A(e_input[23]), .B(g_input[3]), .Z(\mult_23/ab[3][23] ) );
  AND U268 ( .A(e_input[22]), .B(g_input[3]), .Z(\mult_23/ab[3][22] ) );
  AND U269 ( .A(e_input[21]), .B(g_input[3]), .Z(\mult_23/ab[3][21] ) );
  AND U270 ( .A(e_input[20]), .B(g_input[3]), .Z(\mult_23/ab[3][20] ) );
  AND U271 ( .A(e_input[1]), .B(g_input[3]), .Z(\mult_23/ab[3][1] ) );
  AND U272 ( .A(e_input[19]), .B(g_input[3]), .Z(\mult_23/ab[3][19] ) );
  AND U273 ( .A(e_input[18]), .B(g_input[3]), .Z(\mult_23/ab[3][18] ) );
  AND U274 ( .A(e_input[17]), .B(g_input[3]), .Z(\mult_23/ab[3][17] ) );
  AND U275 ( .A(e_input[16]), .B(g_input[3]), .Z(\mult_23/ab[3][16] ) );
  AND U276 ( .A(e_input[15]), .B(g_input[3]), .Z(\mult_23/ab[3][15] ) );
  AND U277 ( .A(e_input[14]), .B(g_input[3]), .Z(\mult_23/ab[3][14] ) );
  AND U278 ( .A(e_input[13]), .B(g_input[3]), .Z(\mult_23/ab[3][13] ) );
  AND U279 ( .A(e_input[12]), .B(g_input[3]), .Z(\mult_23/ab[3][12] ) );
  AND U280 ( .A(e_input[11]), .B(g_input[3]), .Z(\mult_23/ab[3][11] ) );
  AND U281 ( .A(e_input[10]), .B(g_input[3]), .Z(\mult_23/ab[3][10] ) );
  AND U282 ( .A(e_input[0]), .B(g_input[3]), .Z(\mult_23/ab[3][0] ) );
  AND U283 ( .A(g_input[31]), .B(e_input[0]), .Z(\mult_23/ab[31][0] ) );
  AND U284 ( .A(e_input[1]), .B(g_input[30]), .Z(\mult_23/ab[30][1] ) );
  AND U285 ( .A(g_input[30]), .B(e_input[0]), .Z(\mult_23/ab[30][0] ) );
  AND U286 ( .A(e_input[9]), .B(g_input[2]), .Z(\mult_23/ab[2][9] ) );
  AND U287 ( .A(e_input[8]), .B(g_input[2]), .Z(\mult_23/ab[2][8] ) );
  AND U288 ( .A(e_input[7]), .B(g_input[2]), .Z(\mult_23/ab[2][7] ) );
  AND U289 ( .A(e_input[6]), .B(g_input[2]), .Z(\mult_23/ab[2][6] ) );
  AND U290 ( .A(e_input[5]), .B(g_input[2]), .Z(\mult_23/ab[2][5] ) );
  AND U291 ( .A(e_input[4]), .B(g_input[2]), .Z(\mult_23/ab[2][4] ) );
  AND U292 ( .A(e_input[3]), .B(g_input[2]), .Z(\mult_23/ab[2][3] ) );
  AND U293 ( .A(e_input[2]), .B(g_input[2]), .Z(\mult_23/ab[2][2] ) );
  AND U294 ( .A(g_input[2]), .B(e_input[29]), .Z(\mult_23/ab[2][29] ) );
  AND U295 ( .A(e_input[28]), .B(g_input[2]), .Z(\mult_23/ab[2][28] ) );
  AND U296 ( .A(e_input[27]), .B(g_input[2]), .Z(\mult_23/ab[2][27] ) );
  AND U297 ( .A(e_input[26]), .B(g_input[2]), .Z(\mult_23/ab[2][26] ) );
  AND U298 ( .A(e_input[25]), .B(g_input[2]), .Z(\mult_23/ab[2][25] ) );
  AND U299 ( .A(e_input[24]), .B(g_input[2]), .Z(\mult_23/ab[2][24] ) );
  AND U300 ( .A(e_input[23]), .B(g_input[2]), .Z(\mult_23/ab[2][23] ) );
  AND U301 ( .A(e_input[22]), .B(g_input[2]), .Z(\mult_23/ab[2][22] ) );
  AND U302 ( .A(e_input[21]), .B(g_input[2]), .Z(\mult_23/ab[2][21] ) );
  AND U303 ( .A(e_input[20]), .B(g_input[2]), .Z(\mult_23/ab[2][20] ) );
  AND U304 ( .A(e_input[1]), .B(g_input[2]), .Z(\mult_23/ab[2][1] ) );
  AND U305 ( .A(e_input[19]), .B(g_input[2]), .Z(\mult_23/ab[2][19] ) );
  AND U306 ( .A(e_input[18]), .B(g_input[2]), .Z(\mult_23/ab[2][18] ) );
  AND U307 ( .A(e_input[17]), .B(g_input[2]), .Z(\mult_23/ab[2][17] ) );
  AND U308 ( .A(e_input[16]), .B(g_input[2]), .Z(\mult_23/ab[2][16] ) );
  AND U309 ( .A(e_input[15]), .B(g_input[2]), .Z(\mult_23/ab[2][15] ) );
  AND U310 ( .A(e_input[14]), .B(g_input[2]), .Z(\mult_23/ab[2][14] ) );
  AND U311 ( .A(e_input[13]), .B(g_input[2]), .Z(\mult_23/ab[2][13] ) );
  AND U312 ( .A(e_input[12]), .B(g_input[2]), .Z(\mult_23/ab[2][12] ) );
  AND U313 ( .A(e_input[11]), .B(g_input[2]), .Z(\mult_23/ab[2][11] ) );
  AND U314 ( .A(e_input[10]), .B(g_input[2]), .Z(\mult_23/ab[2][10] ) );
  AND U315 ( .A(e_input[0]), .B(g_input[2]), .Z(\mult_23/ab[2][0] ) );
  AND U316 ( .A(e_input[2]), .B(g_input[29]), .Z(\mult_23/ab[29][2] ) );
  AND U317 ( .A(e_input[1]), .B(g_input[29]), .Z(\mult_23/ab[29][1] ) );
  AND U318 ( .A(g_input[29]), .B(e_input[0]), .Z(\mult_23/ab[29][0] ) );
  AND U319 ( .A(e_input[3]), .B(g_input[28]), .Z(\mult_23/ab[28][3] ) );
  AND U320 ( .A(e_input[2]), .B(g_input[28]), .Z(\mult_23/ab[28][2] ) );
  AND U321 ( .A(e_input[1]), .B(g_input[28]), .Z(\mult_23/ab[28][1] ) );
  AND U322 ( .A(g_input[28]), .B(e_input[0]), .Z(\mult_23/ab[28][0] ) );
  AND U323 ( .A(e_input[4]), .B(g_input[27]), .Z(\mult_23/ab[27][4] ) );
  AND U324 ( .A(e_input[3]), .B(g_input[27]), .Z(\mult_23/ab[27][3] ) );
  AND U325 ( .A(e_input[2]), .B(g_input[27]), .Z(\mult_23/ab[27][2] ) );
  AND U326 ( .A(e_input[1]), .B(g_input[27]), .Z(\mult_23/ab[27][1] ) );
  AND U327 ( .A(g_input[27]), .B(e_input[0]), .Z(\mult_23/ab[27][0] ) );
  AND U328 ( .A(e_input[5]), .B(g_input[26]), .Z(\mult_23/ab[26][5] ) );
  AND U329 ( .A(e_input[4]), .B(g_input[26]), .Z(\mult_23/ab[26][4] ) );
  AND U330 ( .A(e_input[3]), .B(g_input[26]), .Z(\mult_23/ab[26][3] ) );
  AND U331 ( .A(e_input[2]), .B(g_input[26]), .Z(\mult_23/ab[26][2] ) );
  AND U332 ( .A(e_input[1]), .B(g_input[26]), .Z(\mult_23/ab[26][1] ) );
  AND U333 ( .A(g_input[26]), .B(e_input[0]), .Z(\mult_23/ab[26][0] ) );
  AND U334 ( .A(e_input[6]), .B(g_input[25]), .Z(\mult_23/ab[25][6] ) );
  AND U335 ( .A(e_input[5]), .B(g_input[25]), .Z(\mult_23/ab[25][5] ) );
  AND U336 ( .A(e_input[4]), .B(g_input[25]), .Z(\mult_23/ab[25][4] ) );
  AND U337 ( .A(e_input[3]), .B(g_input[25]), .Z(\mult_23/ab[25][3] ) );
  AND U338 ( .A(e_input[2]), .B(g_input[25]), .Z(\mult_23/ab[25][2] ) );
  AND U339 ( .A(e_input[1]), .B(g_input[25]), .Z(\mult_23/ab[25][1] ) );
  AND U340 ( .A(g_input[25]), .B(e_input[0]), .Z(\mult_23/ab[25][0] ) );
  AND U341 ( .A(e_input[7]), .B(g_input[24]), .Z(\mult_23/ab[24][7] ) );
  AND U342 ( .A(e_input[6]), .B(g_input[24]), .Z(\mult_23/ab[24][6] ) );
  AND U343 ( .A(e_input[5]), .B(g_input[24]), .Z(\mult_23/ab[24][5] ) );
  AND U344 ( .A(e_input[4]), .B(g_input[24]), .Z(\mult_23/ab[24][4] ) );
  AND U345 ( .A(e_input[3]), .B(g_input[24]), .Z(\mult_23/ab[24][3] ) );
  AND U346 ( .A(e_input[2]), .B(g_input[24]), .Z(\mult_23/ab[24][2] ) );
  AND U347 ( .A(e_input[1]), .B(g_input[24]), .Z(\mult_23/ab[24][1] ) );
  AND U348 ( .A(g_input[24]), .B(e_input[0]), .Z(\mult_23/ab[24][0] ) );
  AND U349 ( .A(e_input[8]), .B(g_input[23]), .Z(\mult_23/ab[23][8] ) );
  AND U350 ( .A(e_input[7]), .B(g_input[23]), .Z(\mult_23/ab[23][7] ) );
  AND U351 ( .A(e_input[6]), .B(g_input[23]), .Z(\mult_23/ab[23][6] ) );
  AND U352 ( .A(e_input[5]), .B(g_input[23]), .Z(\mult_23/ab[23][5] ) );
  AND U353 ( .A(e_input[4]), .B(g_input[23]), .Z(\mult_23/ab[23][4] ) );
  AND U354 ( .A(e_input[3]), .B(g_input[23]), .Z(\mult_23/ab[23][3] ) );
  AND U355 ( .A(e_input[2]), .B(g_input[23]), .Z(\mult_23/ab[23][2] ) );
  AND U356 ( .A(e_input[1]), .B(g_input[23]), .Z(\mult_23/ab[23][1] ) );
  AND U357 ( .A(g_input[23]), .B(e_input[0]), .Z(\mult_23/ab[23][0] ) );
  AND U358 ( .A(e_input[9]), .B(g_input[22]), .Z(\mult_23/ab[22][9] ) );
  AND U359 ( .A(e_input[8]), .B(g_input[22]), .Z(\mult_23/ab[22][8] ) );
  AND U360 ( .A(e_input[7]), .B(g_input[22]), .Z(\mult_23/ab[22][7] ) );
  AND U361 ( .A(e_input[6]), .B(g_input[22]), .Z(\mult_23/ab[22][6] ) );
  AND U362 ( .A(e_input[5]), .B(g_input[22]), .Z(\mult_23/ab[22][5] ) );
  AND U363 ( .A(e_input[4]), .B(g_input[22]), .Z(\mult_23/ab[22][4] ) );
  AND U364 ( .A(e_input[3]), .B(g_input[22]), .Z(\mult_23/ab[22][3] ) );
  AND U365 ( .A(e_input[2]), .B(g_input[22]), .Z(\mult_23/ab[22][2] ) );
  AND U366 ( .A(e_input[1]), .B(g_input[22]), .Z(\mult_23/ab[22][1] ) );
  AND U367 ( .A(g_input[22]), .B(e_input[0]), .Z(\mult_23/ab[22][0] ) );
  AND U368 ( .A(e_input[9]), .B(g_input[21]), .Z(\mult_23/ab[21][9] ) );
  AND U369 ( .A(e_input[8]), .B(g_input[21]), .Z(\mult_23/ab[21][8] ) );
  AND U370 ( .A(e_input[7]), .B(g_input[21]), .Z(\mult_23/ab[21][7] ) );
  AND U371 ( .A(e_input[6]), .B(g_input[21]), .Z(\mult_23/ab[21][6] ) );
  AND U372 ( .A(e_input[5]), .B(g_input[21]), .Z(\mult_23/ab[21][5] ) );
  AND U373 ( .A(e_input[4]), .B(g_input[21]), .Z(\mult_23/ab[21][4] ) );
  AND U374 ( .A(e_input[3]), .B(g_input[21]), .Z(\mult_23/ab[21][3] ) );
  AND U375 ( .A(e_input[2]), .B(g_input[21]), .Z(\mult_23/ab[21][2] ) );
  AND U376 ( .A(e_input[1]), .B(g_input[21]), .Z(\mult_23/ab[21][1] ) );
  AND U377 ( .A(e_input[10]), .B(g_input[21]), .Z(\mult_23/ab[21][10] ) );
  AND U378 ( .A(g_input[21]), .B(e_input[0]), .Z(\mult_23/ab[21][0] ) );
  AND U379 ( .A(e_input[9]), .B(g_input[20]), .Z(\mult_23/ab[20][9] ) );
  AND U380 ( .A(e_input[8]), .B(g_input[20]), .Z(\mult_23/ab[20][8] ) );
  AND U381 ( .A(e_input[7]), .B(g_input[20]), .Z(\mult_23/ab[20][7] ) );
  AND U382 ( .A(e_input[6]), .B(g_input[20]), .Z(\mult_23/ab[20][6] ) );
  AND U383 ( .A(e_input[5]), .B(g_input[20]), .Z(\mult_23/ab[20][5] ) );
  AND U384 ( .A(e_input[4]), .B(g_input[20]), .Z(\mult_23/ab[20][4] ) );
  AND U385 ( .A(e_input[3]), .B(g_input[20]), .Z(\mult_23/ab[20][3] ) );
  AND U386 ( .A(e_input[2]), .B(g_input[20]), .Z(\mult_23/ab[20][2] ) );
  AND U387 ( .A(e_input[1]), .B(g_input[20]), .Z(\mult_23/ab[20][1] ) );
  AND U388 ( .A(e_input[11]), .B(g_input[20]), .Z(\mult_23/ab[20][11] ) );
  AND U389 ( .A(e_input[10]), .B(g_input[20]), .Z(\mult_23/ab[20][10] ) );
  AND U390 ( .A(g_input[20]), .B(e_input[0]), .Z(\mult_23/ab[20][0] ) );
  AND U391 ( .A(e_input[9]), .B(g_input[1]), .Z(\mult_23/ab[1][9] ) );
  AND U392 ( .A(e_input[8]), .B(g_input[1]), .Z(\mult_23/ab[1][8] ) );
  AND U393 ( .A(e_input[7]), .B(g_input[1]), .Z(\mult_23/ab[1][7] ) );
  AND U394 ( .A(e_input[6]), .B(g_input[1]), .Z(\mult_23/ab[1][6] ) );
  AND U395 ( .A(e_input[5]), .B(g_input[1]), .Z(\mult_23/ab[1][5] ) );
  AND U396 ( .A(e_input[4]), .B(g_input[1]), .Z(\mult_23/ab[1][4] ) );
  AND U397 ( .A(e_input[3]), .B(g_input[1]), .Z(\mult_23/ab[1][3] ) );
  AND U398 ( .A(g_input[1]), .B(e_input[30]), .Z(\mult_23/ab[1][30] ) );
  AND U399 ( .A(e_input[2]), .B(g_input[1]), .Z(\mult_23/ab[1][2] ) );
  AND U400 ( .A(e_input[29]), .B(g_input[1]), .Z(\mult_23/ab[1][29] ) );
  AND U401 ( .A(e_input[28]), .B(g_input[1]), .Z(\mult_23/ab[1][28] ) );
  AND U402 ( .A(e_input[27]), .B(g_input[1]), .Z(\mult_23/ab[1][27] ) );
  AND U403 ( .A(e_input[26]), .B(g_input[1]), .Z(\mult_23/ab[1][26] ) );
  AND U404 ( .A(e_input[25]), .B(g_input[1]), .Z(\mult_23/ab[1][25] ) );
  AND U405 ( .A(e_input[24]), .B(g_input[1]), .Z(\mult_23/ab[1][24] ) );
  AND U406 ( .A(e_input[23]), .B(g_input[1]), .Z(\mult_23/ab[1][23] ) );
  AND U407 ( .A(e_input[22]), .B(g_input[1]), .Z(\mult_23/ab[1][22] ) );
  AND U408 ( .A(e_input[21]), .B(g_input[1]), .Z(\mult_23/ab[1][21] ) );
  AND U409 ( .A(e_input[20]), .B(g_input[1]), .Z(\mult_23/ab[1][20] ) );
  AND U410 ( .A(e_input[1]), .B(g_input[1]), .Z(\mult_23/ab[1][1] ) );
  AND U411 ( .A(e_input[19]), .B(g_input[1]), .Z(\mult_23/ab[1][19] ) );
  AND U412 ( .A(e_input[18]), .B(g_input[1]), .Z(\mult_23/ab[1][18] ) );
  AND U413 ( .A(e_input[17]), .B(g_input[1]), .Z(\mult_23/ab[1][17] ) );
  AND U414 ( .A(e_input[16]), .B(g_input[1]), .Z(\mult_23/ab[1][16] ) );
  AND U415 ( .A(e_input[15]), .B(g_input[1]), .Z(\mult_23/ab[1][15] ) );
  AND U416 ( .A(e_input[14]), .B(g_input[1]), .Z(\mult_23/ab[1][14] ) );
  AND U417 ( .A(e_input[13]), .B(g_input[1]), .Z(\mult_23/ab[1][13] ) );
  AND U418 ( .A(e_input[12]), .B(g_input[1]), .Z(\mult_23/ab[1][12] ) );
  AND U419 ( .A(e_input[11]), .B(g_input[1]), .Z(\mult_23/ab[1][11] ) );
  AND U420 ( .A(e_input[10]), .B(g_input[1]), .Z(\mult_23/ab[1][10] ) );
  AND U421 ( .A(e_input[0]), .B(g_input[1]), .Z(\mult_23/ab[1][0] ) );
  AND U422 ( .A(e_input[9]), .B(g_input[19]), .Z(\mult_23/ab[19][9] ) );
  AND U423 ( .A(e_input[8]), .B(g_input[19]), .Z(\mult_23/ab[19][8] ) );
  AND U424 ( .A(e_input[7]), .B(g_input[19]), .Z(\mult_23/ab[19][7] ) );
  AND U425 ( .A(e_input[6]), .B(g_input[19]), .Z(\mult_23/ab[19][6] ) );
  AND U426 ( .A(e_input[5]), .B(g_input[19]), .Z(\mult_23/ab[19][5] ) );
  AND U427 ( .A(e_input[4]), .B(g_input[19]), .Z(\mult_23/ab[19][4] ) );
  AND U428 ( .A(e_input[3]), .B(g_input[19]), .Z(\mult_23/ab[19][3] ) );
  AND U429 ( .A(e_input[2]), .B(g_input[19]), .Z(\mult_23/ab[19][2] ) );
  AND U430 ( .A(e_input[1]), .B(g_input[19]), .Z(\mult_23/ab[19][1] ) );
  AND U431 ( .A(e_input[12]), .B(g_input[19]), .Z(\mult_23/ab[19][12] ) );
  AND U432 ( .A(e_input[11]), .B(g_input[19]), .Z(\mult_23/ab[19][11] ) );
  AND U433 ( .A(e_input[10]), .B(g_input[19]), .Z(\mult_23/ab[19][10] ) );
  AND U434 ( .A(g_input[19]), .B(e_input[0]), .Z(\mult_23/ab[19][0] ) );
  AND U435 ( .A(e_input[9]), .B(g_input[18]), .Z(\mult_23/ab[18][9] ) );
  AND U436 ( .A(e_input[8]), .B(g_input[18]), .Z(\mult_23/ab[18][8] ) );
  AND U437 ( .A(e_input[7]), .B(g_input[18]), .Z(\mult_23/ab[18][7] ) );
  AND U438 ( .A(e_input[6]), .B(g_input[18]), .Z(\mult_23/ab[18][6] ) );
  AND U439 ( .A(e_input[5]), .B(g_input[18]), .Z(\mult_23/ab[18][5] ) );
  AND U440 ( .A(e_input[4]), .B(g_input[18]), .Z(\mult_23/ab[18][4] ) );
  AND U441 ( .A(e_input[3]), .B(g_input[18]), .Z(\mult_23/ab[18][3] ) );
  AND U442 ( .A(e_input[2]), .B(g_input[18]), .Z(\mult_23/ab[18][2] ) );
  AND U443 ( .A(e_input[1]), .B(g_input[18]), .Z(\mult_23/ab[18][1] ) );
  AND U444 ( .A(e_input[13]), .B(g_input[18]), .Z(\mult_23/ab[18][13] ) );
  AND U445 ( .A(e_input[12]), .B(g_input[18]), .Z(\mult_23/ab[18][12] ) );
  AND U446 ( .A(e_input[11]), .B(g_input[18]), .Z(\mult_23/ab[18][11] ) );
  AND U447 ( .A(e_input[10]), .B(g_input[18]), .Z(\mult_23/ab[18][10] ) );
  AND U448 ( .A(g_input[18]), .B(e_input[0]), .Z(\mult_23/ab[18][0] ) );
  AND U449 ( .A(e_input[9]), .B(g_input[17]), .Z(\mult_23/ab[17][9] ) );
  AND U450 ( .A(e_input[8]), .B(g_input[17]), .Z(\mult_23/ab[17][8] ) );
  AND U451 ( .A(e_input[7]), .B(g_input[17]), .Z(\mult_23/ab[17][7] ) );
  AND U452 ( .A(e_input[6]), .B(g_input[17]), .Z(\mult_23/ab[17][6] ) );
  AND U453 ( .A(e_input[5]), .B(g_input[17]), .Z(\mult_23/ab[17][5] ) );
  AND U454 ( .A(e_input[4]), .B(g_input[17]), .Z(\mult_23/ab[17][4] ) );
  AND U455 ( .A(e_input[3]), .B(g_input[17]), .Z(\mult_23/ab[17][3] ) );
  AND U456 ( .A(e_input[2]), .B(g_input[17]), .Z(\mult_23/ab[17][2] ) );
  AND U457 ( .A(e_input[1]), .B(g_input[17]), .Z(\mult_23/ab[17][1] ) );
  AND U458 ( .A(e_input[14]), .B(g_input[17]), .Z(\mult_23/ab[17][14] ) );
  AND U459 ( .A(e_input[13]), .B(g_input[17]), .Z(\mult_23/ab[17][13] ) );
  AND U460 ( .A(e_input[12]), .B(g_input[17]), .Z(\mult_23/ab[17][12] ) );
  AND U461 ( .A(e_input[11]), .B(g_input[17]), .Z(\mult_23/ab[17][11] ) );
  AND U462 ( .A(e_input[10]), .B(g_input[17]), .Z(\mult_23/ab[17][10] ) );
  AND U463 ( .A(g_input[17]), .B(e_input[0]), .Z(\mult_23/ab[17][0] ) );
  AND U464 ( .A(e_input[9]), .B(g_input[16]), .Z(\mult_23/ab[16][9] ) );
  AND U465 ( .A(e_input[8]), .B(g_input[16]), .Z(\mult_23/ab[16][8] ) );
  AND U466 ( .A(e_input[7]), .B(g_input[16]), .Z(\mult_23/ab[16][7] ) );
  AND U467 ( .A(e_input[6]), .B(g_input[16]), .Z(\mult_23/ab[16][6] ) );
  AND U468 ( .A(e_input[5]), .B(g_input[16]), .Z(\mult_23/ab[16][5] ) );
  AND U469 ( .A(e_input[4]), .B(g_input[16]), .Z(\mult_23/ab[16][4] ) );
  AND U470 ( .A(e_input[3]), .B(g_input[16]), .Z(\mult_23/ab[16][3] ) );
  AND U471 ( .A(e_input[2]), .B(g_input[16]), .Z(\mult_23/ab[16][2] ) );
  AND U472 ( .A(e_input[1]), .B(g_input[16]), .Z(\mult_23/ab[16][1] ) );
  AND U473 ( .A(e_input[15]), .B(g_input[16]), .Z(\mult_23/ab[16][15] ) );
  AND U474 ( .A(e_input[14]), .B(g_input[16]), .Z(\mult_23/ab[16][14] ) );
  AND U475 ( .A(e_input[13]), .B(g_input[16]), .Z(\mult_23/ab[16][13] ) );
  AND U476 ( .A(e_input[12]), .B(g_input[16]), .Z(\mult_23/ab[16][12] ) );
  AND U477 ( .A(e_input[11]), .B(g_input[16]), .Z(\mult_23/ab[16][11] ) );
  AND U478 ( .A(e_input[10]), .B(g_input[16]), .Z(\mult_23/ab[16][10] ) );
  AND U479 ( .A(g_input[16]), .B(e_input[0]), .Z(\mult_23/ab[16][0] ) );
  AND U480 ( .A(e_input[9]), .B(g_input[15]), .Z(\mult_23/ab[15][9] ) );
  AND U481 ( .A(e_input[8]), .B(g_input[15]), .Z(\mult_23/ab[15][8] ) );
  AND U482 ( .A(e_input[7]), .B(g_input[15]), .Z(\mult_23/ab[15][7] ) );
  AND U483 ( .A(e_input[6]), .B(g_input[15]), .Z(\mult_23/ab[15][6] ) );
  AND U484 ( .A(e_input[5]), .B(g_input[15]), .Z(\mult_23/ab[15][5] ) );
  AND U485 ( .A(e_input[4]), .B(g_input[15]), .Z(\mult_23/ab[15][4] ) );
  AND U486 ( .A(e_input[3]), .B(g_input[15]), .Z(\mult_23/ab[15][3] ) );
  AND U487 ( .A(e_input[2]), .B(g_input[15]), .Z(\mult_23/ab[15][2] ) );
  AND U488 ( .A(e_input[1]), .B(g_input[15]), .Z(\mult_23/ab[15][1] ) );
  AND U489 ( .A(e_input[16]), .B(g_input[15]), .Z(\mult_23/ab[15][16] ) );
  AND U490 ( .A(e_input[15]), .B(g_input[15]), .Z(\mult_23/ab[15][15] ) );
  AND U491 ( .A(e_input[14]), .B(g_input[15]), .Z(\mult_23/ab[15][14] ) );
  AND U492 ( .A(e_input[13]), .B(g_input[15]), .Z(\mult_23/ab[15][13] ) );
  AND U493 ( .A(e_input[12]), .B(g_input[15]), .Z(\mult_23/ab[15][12] ) );
  AND U494 ( .A(e_input[11]), .B(g_input[15]), .Z(\mult_23/ab[15][11] ) );
  AND U495 ( .A(e_input[10]), .B(g_input[15]), .Z(\mult_23/ab[15][10] ) );
  AND U496 ( .A(g_input[15]), .B(e_input[0]), .Z(\mult_23/ab[15][0] ) );
  AND U497 ( .A(e_input[9]), .B(g_input[14]), .Z(\mult_23/ab[14][9] ) );
  AND U498 ( .A(e_input[8]), .B(g_input[14]), .Z(\mult_23/ab[14][8] ) );
  AND U499 ( .A(e_input[7]), .B(g_input[14]), .Z(\mult_23/ab[14][7] ) );
  AND U500 ( .A(e_input[6]), .B(g_input[14]), .Z(\mult_23/ab[14][6] ) );
  AND U501 ( .A(e_input[5]), .B(g_input[14]), .Z(\mult_23/ab[14][5] ) );
  AND U502 ( .A(e_input[4]), .B(g_input[14]), .Z(\mult_23/ab[14][4] ) );
  AND U503 ( .A(e_input[3]), .B(g_input[14]), .Z(\mult_23/ab[14][3] ) );
  AND U504 ( .A(e_input[2]), .B(g_input[14]), .Z(\mult_23/ab[14][2] ) );
  AND U505 ( .A(e_input[1]), .B(g_input[14]), .Z(\mult_23/ab[14][1] ) );
  AND U506 ( .A(e_input[17]), .B(g_input[14]), .Z(\mult_23/ab[14][17] ) );
  AND U507 ( .A(e_input[16]), .B(g_input[14]), .Z(\mult_23/ab[14][16] ) );
  AND U508 ( .A(e_input[15]), .B(g_input[14]), .Z(\mult_23/ab[14][15] ) );
  AND U509 ( .A(e_input[14]), .B(g_input[14]), .Z(\mult_23/ab[14][14] ) );
  AND U510 ( .A(e_input[13]), .B(g_input[14]), .Z(\mult_23/ab[14][13] ) );
  AND U511 ( .A(e_input[12]), .B(g_input[14]), .Z(\mult_23/ab[14][12] ) );
  AND U512 ( .A(e_input[11]), .B(g_input[14]), .Z(\mult_23/ab[14][11] ) );
  AND U513 ( .A(e_input[10]), .B(g_input[14]), .Z(\mult_23/ab[14][10] ) );
  AND U514 ( .A(g_input[14]), .B(e_input[0]), .Z(\mult_23/ab[14][0] ) );
  AND U515 ( .A(e_input[9]), .B(g_input[13]), .Z(\mult_23/ab[13][9] ) );
  AND U516 ( .A(e_input[8]), .B(g_input[13]), .Z(\mult_23/ab[13][8] ) );
  AND U517 ( .A(e_input[7]), .B(g_input[13]), .Z(\mult_23/ab[13][7] ) );
  AND U518 ( .A(e_input[6]), .B(g_input[13]), .Z(\mult_23/ab[13][6] ) );
  AND U519 ( .A(e_input[5]), .B(g_input[13]), .Z(\mult_23/ab[13][5] ) );
  AND U520 ( .A(e_input[4]), .B(g_input[13]), .Z(\mult_23/ab[13][4] ) );
  AND U521 ( .A(e_input[3]), .B(g_input[13]), .Z(\mult_23/ab[13][3] ) );
  AND U522 ( .A(e_input[2]), .B(g_input[13]), .Z(\mult_23/ab[13][2] ) );
  AND U523 ( .A(e_input[1]), .B(g_input[13]), .Z(\mult_23/ab[13][1] ) );
  AND U524 ( .A(e_input[18]), .B(g_input[13]), .Z(\mult_23/ab[13][18] ) );
  AND U525 ( .A(e_input[17]), .B(g_input[13]), .Z(\mult_23/ab[13][17] ) );
  AND U526 ( .A(e_input[16]), .B(g_input[13]), .Z(\mult_23/ab[13][16] ) );
  AND U527 ( .A(e_input[15]), .B(g_input[13]), .Z(\mult_23/ab[13][15] ) );
  AND U528 ( .A(e_input[14]), .B(g_input[13]), .Z(\mult_23/ab[13][14] ) );
  AND U529 ( .A(e_input[13]), .B(g_input[13]), .Z(\mult_23/ab[13][13] ) );
  AND U530 ( .A(e_input[12]), .B(g_input[13]), .Z(\mult_23/ab[13][12] ) );
  AND U531 ( .A(e_input[11]), .B(g_input[13]), .Z(\mult_23/ab[13][11] ) );
  AND U532 ( .A(e_input[10]), .B(g_input[13]), .Z(\mult_23/ab[13][10] ) );
  AND U533 ( .A(g_input[13]), .B(e_input[0]), .Z(\mult_23/ab[13][0] ) );
  AND U534 ( .A(e_input[9]), .B(g_input[12]), .Z(\mult_23/ab[12][9] ) );
  AND U535 ( .A(e_input[8]), .B(g_input[12]), .Z(\mult_23/ab[12][8] ) );
  AND U536 ( .A(e_input[7]), .B(g_input[12]), .Z(\mult_23/ab[12][7] ) );
  AND U537 ( .A(e_input[6]), .B(g_input[12]), .Z(\mult_23/ab[12][6] ) );
  AND U538 ( .A(e_input[5]), .B(g_input[12]), .Z(\mult_23/ab[12][5] ) );
  AND U539 ( .A(e_input[4]), .B(g_input[12]), .Z(\mult_23/ab[12][4] ) );
  AND U540 ( .A(e_input[3]), .B(g_input[12]), .Z(\mult_23/ab[12][3] ) );
  AND U541 ( .A(e_input[2]), .B(g_input[12]), .Z(\mult_23/ab[12][2] ) );
  AND U542 ( .A(e_input[1]), .B(g_input[12]), .Z(\mult_23/ab[12][1] ) );
  AND U543 ( .A(e_input[19]), .B(g_input[12]), .Z(\mult_23/ab[12][19] ) );
  AND U544 ( .A(e_input[18]), .B(g_input[12]), .Z(\mult_23/ab[12][18] ) );
  AND U545 ( .A(e_input[17]), .B(g_input[12]), .Z(\mult_23/ab[12][17] ) );
  AND U546 ( .A(e_input[16]), .B(g_input[12]), .Z(\mult_23/ab[12][16] ) );
  AND U547 ( .A(e_input[15]), .B(g_input[12]), .Z(\mult_23/ab[12][15] ) );
  AND U548 ( .A(e_input[14]), .B(g_input[12]), .Z(\mult_23/ab[12][14] ) );
  AND U549 ( .A(e_input[13]), .B(g_input[12]), .Z(\mult_23/ab[12][13] ) );
  AND U550 ( .A(e_input[12]), .B(g_input[12]), .Z(\mult_23/ab[12][12] ) );
  AND U551 ( .A(e_input[11]), .B(g_input[12]), .Z(\mult_23/ab[12][11] ) );
  AND U552 ( .A(e_input[10]), .B(g_input[12]), .Z(\mult_23/ab[12][10] ) );
  AND U553 ( .A(g_input[12]), .B(e_input[0]), .Z(\mult_23/ab[12][0] ) );
  AND U554 ( .A(e_input[9]), .B(g_input[11]), .Z(\mult_23/ab[11][9] ) );
  AND U555 ( .A(e_input[8]), .B(g_input[11]), .Z(\mult_23/ab[11][8] ) );
  AND U556 ( .A(e_input[7]), .B(g_input[11]), .Z(\mult_23/ab[11][7] ) );
  AND U557 ( .A(e_input[6]), .B(g_input[11]), .Z(\mult_23/ab[11][6] ) );
  AND U558 ( .A(e_input[5]), .B(g_input[11]), .Z(\mult_23/ab[11][5] ) );
  AND U559 ( .A(e_input[4]), .B(g_input[11]), .Z(\mult_23/ab[11][4] ) );
  AND U560 ( .A(e_input[3]), .B(g_input[11]), .Z(\mult_23/ab[11][3] ) );
  AND U561 ( .A(e_input[2]), .B(g_input[11]), .Z(\mult_23/ab[11][2] ) );
  AND U562 ( .A(e_input[20]), .B(g_input[11]), .Z(\mult_23/ab[11][20] ) );
  AND U563 ( .A(e_input[1]), .B(g_input[11]), .Z(\mult_23/ab[11][1] ) );
  AND U564 ( .A(e_input[19]), .B(g_input[11]), .Z(\mult_23/ab[11][19] ) );
  AND U565 ( .A(e_input[18]), .B(g_input[11]), .Z(\mult_23/ab[11][18] ) );
  AND U566 ( .A(e_input[17]), .B(g_input[11]), .Z(\mult_23/ab[11][17] ) );
  AND U567 ( .A(e_input[16]), .B(g_input[11]), .Z(\mult_23/ab[11][16] ) );
  AND U568 ( .A(e_input[15]), .B(g_input[11]), .Z(\mult_23/ab[11][15] ) );
  AND U569 ( .A(e_input[14]), .B(g_input[11]), .Z(\mult_23/ab[11][14] ) );
  AND U570 ( .A(e_input[13]), .B(g_input[11]), .Z(\mult_23/ab[11][13] ) );
  AND U571 ( .A(e_input[12]), .B(g_input[11]), .Z(\mult_23/ab[11][12] ) );
  AND U572 ( .A(e_input[11]), .B(g_input[11]), .Z(\mult_23/ab[11][11] ) );
  AND U573 ( .A(e_input[10]), .B(g_input[11]), .Z(\mult_23/ab[11][10] ) );
  AND U574 ( .A(g_input[11]), .B(e_input[0]), .Z(\mult_23/ab[11][0] ) );
  AND U575 ( .A(e_input[9]), .B(g_input[10]), .Z(\mult_23/ab[10][9] ) );
  AND U576 ( .A(e_input[8]), .B(g_input[10]), .Z(\mult_23/ab[10][8] ) );
  AND U577 ( .A(e_input[7]), .B(g_input[10]), .Z(\mult_23/ab[10][7] ) );
  AND U578 ( .A(e_input[6]), .B(g_input[10]), .Z(\mult_23/ab[10][6] ) );
  AND U579 ( .A(e_input[5]), .B(g_input[10]), .Z(\mult_23/ab[10][5] ) );
  AND U580 ( .A(e_input[4]), .B(g_input[10]), .Z(\mult_23/ab[10][4] ) );
  AND U581 ( .A(e_input[3]), .B(g_input[10]), .Z(\mult_23/ab[10][3] ) );
  AND U582 ( .A(e_input[2]), .B(g_input[10]), .Z(\mult_23/ab[10][2] ) );
  AND U583 ( .A(e_input[21]), .B(g_input[10]), .Z(\mult_23/ab[10][21] ) );
  AND U584 ( .A(e_input[20]), .B(g_input[10]), .Z(\mult_23/ab[10][20] ) );
  AND U585 ( .A(e_input[1]), .B(g_input[10]), .Z(\mult_23/ab[10][1] ) );
  AND U586 ( .A(e_input[19]), .B(g_input[10]), .Z(\mult_23/ab[10][19] ) );
  AND U587 ( .A(e_input[18]), .B(g_input[10]), .Z(\mult_23/ab[10][18] ) );
  AND U588 ( .A(e_input[17]), .B(g_input[10]), .Z(\mult_23/ab[10][17] ) );
  AND U589 ( .A(e_input[16]), .B(g_input[10]), .Z(\mult_23/ab[10][16] ) );
  AND U590 ( .A(e_input[15]), .B(g_input[10]), .Z(\mult_23/ab[10][15] ) );
  AND U591 ( .A(e_input[14]), .B(g_input[10]), .Z(\mult_23/ab[10][14] ) );
  AND U592 ( .A(e_input[13]), .B(g_input[10]), .Z(\mult_23/ab[10][13] ) );
  AND U593 ( .A(e_input[12]), .B(g_input[10]), .Z(\mult_23/ab[10][12] ) );
  AND U594 ( .A(e_input[11]), .B(g_input[10]), .Z(\mult_23/ab[10][11] ) );
  AND U595 ( .A(e_input[10]), .B(g_input[10]), .Z(\mult_23/ab[10][10] ) );
  AND U596 ( .A(g_input[10]), .B(e_input[0]), .Z(\mult_23/ab[10][0] ) );
  AND U597 ( .A(g_input[0]), .B(e_input[9]), .Z(\mult_23/ab[0][9] ) );
  AND U598 ( .A(g_input[0]), .B(e_input[8]), .Z(\mult_23/ab[0][8] ) );
  AND U599 ( .A(g_input[0]), .B(e_input[7]), .Z(\mult_23/ab[0][7] ) );
  AND U600 ( .A(g_input[0]), .B(e_input[6]), .Z(\mult_23/ab[0][6] ) );
  AND U601 ( .A(g_input[0]), .B(e_input[5]), .Z(\mult_23/ab[0][5] ) );
  AND U602 ( .A(g_input[0]), .B(e_input[4]), .Z(\mult_23/ab[0][4] ) );
  AND U603 ( .A(g_input[0]), .B(e_input[3]), .Z(\mult_23/ab[0][3] ) );
  AND U604 ( .A(e_input[31]), .B(g_input[0]), .Z(\mult_23/ab[0][31] ) );
  AND U605 ( .A(e_input[30]), .B(g_input[0]), .Z(\mult_23/ab[0][30] ) );
  AND U606 ( .A(g_input[0]), .B(e_input[2]), .Z(\mult_23/ab[0][2] ) );
  AND U607 ( .A(g_input[0]), .B(e_input[29]), .Z(\mult_23/ab[0][29] ) );
  AND U608 ( .A(g_input[0]), .B(e_input[28]), .Z(\mult_23/ab[0][28] ) );
  AND U609 ( .A(g_input[0]), .B(e_input[27]), .Z(\mult_23/ab[0][27] ) );
  AND U610 ( .A(g_input[0]), .B(e_input[26]), .Z(\mult_23/ab[0][26] ) );
  AND U611 ( .A(g_input[0]), .B(e_input[25]), .Z(\mult_23/ab[0][25] ) );
  AND U612 ( .A(g_input[0]), .B(e_input[24]), .Z(\mult_23/ab[0][24] ) );
  AND U613 ( .A(g_input[0]), .B(e_input[23]), .Z(\mult_23/ab[0][23] ) );
  AND U614 ( .A(g_input[0]), .B(e_input[22]), .Z(\mult_23/ab[0][22] ) );
  AND U615 ( .A(g_input[0]), .B(e_input[21]), .Z(\mult_23/ab[0][21] ) );
  AND U616 ( .A(g_input[0]), .B(e_input[20]), .Z(\mult_23/ab[0][20] ) );
  AND U617 ( .A(g_input[0]), .B(e_input[1]), .Z(\mult_23/ab[0][1] ) );
  AND U618 ( .A(g_input[0]), .B(e_input[19]), .Z(\mult_23/ab[0][19] ) );
  AND U619 ( .A(g_input[0]), .B(e_input[18]), .Z(\mult_23/ab[0][18] ) );
  AND U620 ( .A(g_input[0]), .B(e_input[17]), .Z(\mult_23/ab[0][17] ) );
  AND U621 ( .A(g_input[0]), .B(e_input[16]), .Z(\mult_23/ab[0][16] ) );
  AND U622 ( .A(g_input[0]), .B(e_input[15]), .Z(\mult_23/ab[0][15] ) );
  AND U623 ( .A(g_input[0]), .B(e_input[14]), .Z(\mult_23/ab[0][14] ) );
  AND U624 ( .A(g_input[0]), .B(e_input[13]), .Z(\mult_23/ab[0][13] ) );
  AND U625 ( .A(g_input[0]), .B(e_input[12]), .Z(\mult_23/ab[0][12] ) );
  AND U626 ( .A(g_input[0]), .B(e_input[11]), .Z(\mult_23/ab[0][11] ) );
  AND U627 ( .A(g_input[0]), .B(e_input[10]), .Z(\mult_23/ab[0][10] ) );
endmodule

